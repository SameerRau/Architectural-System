<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>5.71504,-22.9877,112.962,-75.9978</PageViewport>
<gate>
<ID>1</ID>
<type>AE_MUX_4x1</type>
<position>38,-11</position>
<input>
<ID>IN_0</ID>7 </input>
<input>
<ID>IN_1</ID>143 </input>
<input>
<ID>IN_2</ID>135 </input>
<input>
<ID>IN_3</ID>127 </input>
<output>
<ID>OUT</ID>87 </output>
<input>
<ID>SEL_0</ID>94 </input>
<input>
<ID>SEL_1</ID>93 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>2</ID>
<type>AE_MUX_4x1</type>
<position>38,-22</position>
<input>
<ID>IN_0</ID>6 </input>
<input>
<ID>IN_1</ID>144 </input>
<input>
<ID>IN_2</ID>136 </input>
<input>
<ID>IN_3</ID>128 </input>
<output>
<ID>OUT</ID>86 </output>
<input>
<ID>SEL_0</ID>94 </input>
<input>
<ID>SEL_1</ID>93 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>3</ID>
<type>AE_MUX_4x1</type>
<position>38,-33</position>
<input>
<ID>IN_0</ID>5 </input>
<input>
<ID>IN_1</ID>145 </input>
<input>
<ID>IN_2</ID>137 </input>
<input>
<ID>IN_3</ID>129 </input>
<output>
<ID>OUT</ID>85 </output>
<input>
<ID>SEL_0</ID>94 </input>
<input>
<ID>SEL_1</ID>93 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>4</ID>
<type>AE_MUX_4x1</type>
<position>38,-43.5</position>
<input>
<ID>IN_0</ID>4 </input>
<input>
<ID>IN_1</ID>146 </input>
<input>
<ID>IN_2</ID>138 </input>
<input>
<ID>IN_3</ID>130 </input>
<output>
<ID>OUT</ID>80 </output>
<input>
<ID>SEL_0</ID>94 </input>
<input>
<ID>SEL_1</ID>93 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>5</ID>
<type>AE_MUX_4x1</type>
<position>38,-53.5</position>
<input>
<ID>IN_0</ID>3 </input>
<input>
<ID>IN_1</ID>147 </input>
<input>
<ID>IN_2</ID>139 </input>
<input>
<ID>IN_3</ID>131 </input>
<output>
<ID>OUT</ID>79 </output>
<input>
<ID>SEL_0</ID>94 </input>
<input>
<ID>SEL_1</ID>93 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>6</ID>
<type>AE_MUX_4x1</type>
<position>38,-63.5</position>
<input>
<ID>IN_0</ID>2 </input>
<input>
<ID>IN_1</ID>148 </input>
<input>
<ID>IN_2</ID>140 </input>
<input>
<ID>IN_3</ID>133 </input>
<output>
<ID>OUT</ID>78 </output>
<input>
<ID>SEL_0</ID>94 </input>
<input>
<ID>SEL_1</ID>93 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>7</ID>
<type>AE_MUX_4x1</type>
<position>38,-73.5</position>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>149 </input>
<input>
<ID>IN_2</ID>141 </input>
<input>
<ID>IN_3</ID>133 </input>
<output>
<ID>OUT</ID>77 </output>
<input>
<ID>SEL_0</ID>94 </input>
<input>
<ID>SEL_1</ID>93 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>8</ID>
<type>AE_MUX_4x1</type>
<position>48,-11</position>
<input>
<ID>IN_0</ID>7 </input>
<input>
<ID>IN_1</ID>143 </input>
<input>
<ID>IN_2</ID>135 </input>
<input>
<ID>IN_3</ID>127 </input>
<output>
<ID>OUT</ID>91 </output>
<input>
<ID>SEL_0</ID>154 </input>
<input>
<ID>SEL_1</ID>153 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>9</ID>
<type>AE_MUX_4x1</type>
<position>48,-22</position>
<input>
<ID>IN_0</ID>6 </input>
<input>
<ID>IN_1</ID>144 </input>
<input>
<ID>IN_2</ID>136 </input>
<input>
<ID>IN_3</ID>128 </input>
<output>
<ID>OUT</ID>90 </output>
<input>
<ID>SEL_0</ID>154 </input>
<input>
<ID>SEL_1</ID>153 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>10</ID>
<type>AE_MUX_4x1</type>
<position>48,-33</position>
<input>
<ID>IN_0</ID>5 </input>
<input>
<ID>IN_1</ID>145 </input>
<input>
<ID>IN_2</ID>137 </input>
<input>
<ID>IN_3</ID>129 </input>
<output>
<ID>OUT</ID>89 </output>
<input>
<ID>SEL_0</ID>154 </input>
<input>
<ID>SEL_1</ID>153 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>11</ID>
<type>AE_MUX_4x1</type>
<position>48,-43</position>
<input>
<ID>IN_0</ID>4 </input>
<input>
<ID>IN_1</ID>146 </input>
<input>
<ID>IN_2</ID>138 </input>
<input>
<ID>IN_3</ID>130 </input>
<output>
<ID>OUT</ID>84 </output>
<input>
<ID>SEL_0</ID>154 </input>
<input>
<ID>SEL_1</ID>153 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>12</ID>
<type>AE_MUX_4x1</type>
<position>48,-53.5</position>
<input>
<ID>IN_0</ID>3 </input>
<input>
<ID>IN_1</ID>147 </input>
<input>
<ID>IN_2</ID>139 </input>
<input>
<ID>IN_3</ID>131 </input>
<output>
<ID>OUT</ID>83 </output>
<input>
<ID>SEL_0</ID>154 </input>
<input>
<ID>SEL_1</ID>153 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>13</ID>
<type>AE_MUX_4x1</type>
<position>48,-63.5</position>
<input>
<ID>IN_0</ID>2 </input>
<input>
<ID>IN_1</ID>148 </input>
<input>
<ID>IN_2</ID>140 </input>
<input>
<ID>IN_3</ID>133 </input>
<output>
<ID>OUT</ID>82 </output>
<input>
<ID>SEL_0</ID>154 </input>
<input>
<ID>SEL_1</ID>153 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>14</ID>
<type>AE_MUX_4x1</type>
<position>48,-73.5</position>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>149 </input>
<input>
<ID>IN_2</ID>141 </input>
<input>
<ID>IN_3</ID>133 </input>
<output>
<ID>OUT</ID>81 </output>
<input>
<ID>SEL_0</ID>154 </input>
<input>
<ID>SEL_1</ID>153 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>15</ID>
<type>AE_MUX_4x1</type>
<position>48,-1</position>
<input>
<ID>IN_0</ID>8 </input>
<input>
<ID>IN_1</ID>142 </input>
<input>
<ID>IN_2</ID>134 </input>
<input>
<ID>IN_3</ID>126 </input>
<output>
<ID>OUT</ID>92 </output>
<input>
<ID>SEL_0</ID>154 </input>
<input>
<ID>SEL_1</ID>153 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>16</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>61.5,4.5</position>
<input>
<ID>ENABLE_0</ID>9 </input>
<input>
<ID>IN_0</ID>81 </input>
<input>
<ID>IN_1</ID>82 </input>
<input>
<ID>IN_2</ID>83 </input>
<input>
<ID>IN_3</ID>84 </input>
<input>
<ID>IN_4</ID>89 </input>
<input>
<ID>IN_5</ID>90 </input>
<input>
<ID>IN_6</ID>91 </input>
<input>
<ID>IN_7</ID>92 </input>
<output>
<ID>OUT_0</ID>29 </output>
<output>
<ID>OUT_1</ID>30 </output>
<output>
<ID>OUT_2</ID>31 </output>
<output>
<ID>OUT_3</ID>32 </output>
<output>
<ID>OUT_4</ID>33 </output>
<output>
<ID>OUT_5</ID>34 </output>
<output>
<ID>OUT_6</ID>35 </output>
<output>
<ID>OUT_7</ID>36 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>17</ID>
<type>BI_TRI_STATE_4BIT</type>
<position>47.5,26.5</position>
<input>
<ID>ENABLE_0</ID>152 </input>
<input>
<ID>IN_2</ID>93 </input>
<input>
<ID>IN_3</ID>151 </input>
<output>
<ID>OUT_2</ID>153 </output>
<output>
<ID>OUT_3</ID>154 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>18</ID>
<type>AE_SMALL_INVERTER</type>
<position>53,26.5</position>
<input>
<ID>IN_0</ID>9 </input>
<output>
<ID>OUT_0</ID>152 </output>
<gparam>angle 180</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>19</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>-26,-37</position>
<input>
<ID>ENABLE_0</ID>70 </input>
<input>
<ID>IN_0</ID>103 </input>
<input>
<ID>IN_1</ID>19 </input>
<input>
<ID>IN_2</ID>20 </input>
<input>
<ID>IN_3</ID>21 </input>
<input>
<ID>IN_4</ID>22 </input>
<input>
<ID>IN_5</ID>23 </input>
<input>
<ID>IN_6</ID>24 </input>
<input>
<ID>IN_7</ID>25 </input>
<output>
<ID>OUT_0</ID>15 </output>
<output>
<ID>OUT_1</ID>16 </output>
<output>
<ID>OUT_2</ID>17 </output>
<output>
<ID>OUT_3</ID>18 </output>
<output>
<ID>OUT_4</ID>26 </output>
<output>
<ID>OUT_5</ID>27 </output>
<output>
<ID>OUT_6</ID>28 </output>
<output>
<ID>OUT_7</ID>37 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>20</ID>
<type>BI_TRI_STATE_4BIT</type>
<position>41.5,26.5</position>
<input>
<ID>ENABLE_0</ID>9 </input>
<input>
<ID>IN_2</ID>124 </input>
<input>
<ID>IN_3</ID>125 </input>
<output>
<ID>OUT_2</ID>153 </output>
<output>
<ID>OUT_3</ID>154 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>21</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>-26,-25.5</position>
<input>
<ID>ENABLE_0</ID>10 </input>
<input>
<ID>IN_0</ID>29 </input>
<input>
<ID>IN_1</ID>30 </input>
<input>
<ID>IN_2</ID>31 </input>
<input>
<ID>IN_3</ID>32 </input>
<input>
<ID>IN_4</ID>33 </input>
<input>
<ID>IN_5</ID>34 </input>
<input>
<ID>IN_6</ID>35 </input>
<input>
<ID>IN_7</ID>36 </input>
<output>
<ID>OUT_0</ID>15 </output>
<output>
<ID>OUT_1</ID>16 </output>
<output>
<ID>OUT_2</ID>17 </output>
<output>
<ID>OUT_3</ID>18 </output>
<output>
<ID>OUT_4</ID>26 </output>
<output>
<ID>OUT_5</ID>27 </output>
<output>
<ID>OUT_6</ID>28 </output>
<output>
<ID>OUT_7</ID>37 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>22</ID>
<type>AE_REGISTER8</type>
<position>15,-26</position>
<input>
<ID>IN_0</ID>53 </input>
<input>
<ID>IN_1</ID>47 </input>
<input>
<ID>IN_2</ID>46 </input>
<input>
<ID>IN_3</ID>50 </input>
<input>
<ID>IN_4</ID>48 </input>
<input>
<ID>IN_5</ID>49 </input>
<input>
<ID>IN_6</ID>51 </input>
<input>
<ID>IN_7</ID>52 </input>
<output>
<ID>OUT_0</ID>141 </output>
<output>
<ID>OUT_1</ID>140 </output>
<output>
<ID>OUT_2</ID>139 </output>
<output>
<ID>OUT_3</ID>138 </output>
<output>
<ID>OUT_4</ID>137 </output>
<output>
<ID>OUT_5</ID>136 </output>
<output>
<ID>OUT_6</ID>135 </output>
<output>
<ID>OUT_7</ID>134 </output>
<input>
<ID>clock</ID>75 </input>
<input>
<ID>load</ID>73 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 3</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>23</ID>
<type>AE_REGISTER8</type>
<position>15,-46.5</position>
<input>
<ID>IN_0</ID>57 </input>
<input>
<ID>IN_1</ID>61 </input>
<input>
<ID>IN_2</ID>58 </input>
<input>
<ID>IN_3</ID>54 </input>
<input>
<ID>IN_4</ID>59 </input>
<input>
<ID>IN_5</ID>55 </input>
<input>
<ID>IN_6</ID>56 </input>
<input>
<ID>IN_7</ID>60 </input>
<output>
<ID>OUT_0</ID>149 </output>
<output>
<ID>OUT_1</ID>148 </output>
<output>
<ID>OUT_2</ID>147 </output>
<output>
<ID>OUT_3</ID>146 </output>
<output>
<ID>OUT_4</ID>145 </output>
<output>
<ID>OUT_5</ID>144 </output>
<output>
<ID>OUT_6</ID>143 </output>
<output>
<ID>OUT_7</ID>142 </output>
<input>
<ID>clock</ID>75 </input>
<input>
<ID>load</ID>72 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 2</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>24</ID>
<type>AE_REGISTER8</type>
<position>15,-65.5</position>
<input>
<ID>IN_0</ID>64 </input>
<input>
<ID>IN_1</ID>63 </input>
<input>
<ID>IN_2</ID>69 </input>
<input>
<ID>IN_3</ID>65 </input>
<input>
<ID>IN_4</ID>66 </input>
<input>
<ID>IN_5</ID>67 </input>
<input>
<ID>IN_6</ID>62 </input>
<input>
<ID>IN_7</ID>68 </input>
<output>
<ID>OUT_0</ID>1 </output>
<output>
<ID>OUT_1</ID>2 </output>
<output>
<ID>OUT_2</ID>3 </output>
<output>
<ID>OUT_3</ID>4 </output>
<output>
<ID>OUT_4</ID>5 </output>
<output>
<ID>OUT_5</ID>6 </output>
<output>
<ID>OUT_6</ID>7 </output>
<output>
<ID>OUT_7</ID>8 </output>
<input>
<ID>clock</ID>75 </input>
<input>
<ID>load</ID>71 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>25</ID>
<type>BA_DECODER_2x4</type>
<position>-15.5,26.5</position>
<input>
<ID>ENABLE</ID>14 </input>
<input>
<ID>IN_0</ID>125 </input>
<input>
<ID>IN_1</ID>124 </input>
<output>
<ID>OUT_0</ID>71 </output>
<output>
<ID>OUT_1</ID>72 </output>
<output>
<ID>OUT_2</ID>73 </output>
<output>
<ID>OUT_3</ID>74 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>26</ID>
<type>AA_LABEL</type>
<position>46.5,42.5</position>
<gparam>LABEL_TEXT Bits 0 - 5 are for the source registers / destination registers / memory address</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>27</ID>
<type>BA_DECODER_2x4</type>
<position>-15.5,21</position>
<input>
<ID>ENABLE</ID>121 </input>
<input>
<ID>IN_0</ID>122 </input>
<input>
<ID>IN_1</ID>123 </input>
<output>
<ID>OUT_0</ID>9 </output>
<output>
<ID>OUT_1</ID>10 </output>
<output>
<ID>OUT_2</ID>11 </output>
<output>
<ID>OUT_3</ID>13 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>28</ID>
<type>AA_LABEL</type>
<position>28,40.5</position>
<gparam>LABEL_TEXT Bits 6 - 7 are for the opcodes</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>29</ID>
<type>AE_SMALL_INVERTER</type>
<position>101,-3</position>
<input>
<ID>IN_0</ID>11 </input>
<output>
<ID>OUT_0</ID>12 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>30</ID>
<type>AA_AND2</type>
<position>102,-8.5</position>
<input>
<ID>IN_0</ID>13 </input>
<input>
<ID>IN_1</ID>12 </input>
<output>
<ID>OUT</ID>112 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>31</ID>
<type>AE_RAM_8x8</type>
<position>-35.5,14</position>
<input>
<ID>ADDRESS_0</ID>94 </input>
<input>
<ID>ADDRESS_1</ID>93 </input>
<input>
<ID>ADDRESS_2</ID>151 </input>
<input>
<ID>ADDRESS_3</ID>93 </input>
<input>
<ID>ADDRESS_4</ID>125 </input>
<input>
<ID>ADDRESS_5</ID>124 </input>
<input>
<ID>ADDRESS_6</ID>122 </input>
<input>
<ID>ADDRESS_7</ID>123 </input>
<input>
<ID>DATA_IN_0</ID>29 </input>
<input>
<ID>DATA_IN_1</ID>30 </input>
<input>
<ID>DATA_IN_2</ID>31 </input>
<input>
<ID>DATA_IN_3</ID>32 </input>
<input>
<ID>DATA_IN_4</ID>33 </input>
<input>
<ID>DATA_IN_5</ID>34 </input>
<input>
<ID>DATA_IN_6</ID>35 </input>
<input>
<ID>DATA_IN_7</ID>36 </input>
<output>
<ID>DATA_OUT_0</ID>29 </output>
<output>
<ID>DATA_OUT_1</ID>30 </output>
<output>
<ID>DATA_OUT_2</ID>31 </output>
<output>
<ID>DATA_OUT_3</ID>32 </output>
<output>
<ID>DATA_OUT_4</ID>33 </output>
<output>
<ID>DATA_OUT_5</ID>34 </output>
<output>
<ID>DATA_OUT_6</ID>35 </output>
<output>
<ID>DATA_OUT_7</ID>36 </output>
<input>
<ID>ENABLE_0</ID>10 </input>
<input>
<ID>write_clock</ID>75 </input>
<input>
<ID>write_enable</ID>9 </input>
<gparam>angle 0.0</gparam>
<lparam>ADDRESS_BITS 8</lparam>
<lparam>DATA_BITS 8</lparam>
<lparam>Address:0 1</lparam></gate>
<gate>
<ID>32</ID>
<type>BE_ROM_8x8</type>
<position>4,40</position>
<input>
<ID>ADDRESS_0</ID>113 </input>
<input>
<ID>ADDRESS_1</ID>114 </input>
<input>
<ID>ADDRESS_2</ID>115 </input>
<input>
<ID>ADDRESS_3</ID>116 </input>
<input>
<ID>ADDRESS_4</ID>117 </input>
<input>
<ID>ADDRESS_5</ID>118 </input>
<input>
<ID>ADDRESS_6</ID>119 </input>
<input>
<ID>ADDRESS_7</ID>120 </input>
<output>
<ID>DATA_OUT_0</ID>94 </output>
<output>
<ID>DATA_OUT_1</ID>93 </output>
<output>
<ID>DATA_OUT_2</ID>151 </output>
<output>
<ID>DATA_OUT_3</ID>93 </output>
<output>
<ID>DATA_OUT_4</ID>125 </output>
<output>
<ID>DATA_OUT_5</ID>124 </output>
<output>
<ID>DATA_OUT_6</ID>122 </output>
<output>
<ID>DATA_OUT_7</ID>123 </output>
<input>
<ID>ENABLE_0</ID>121 </input>
<gparam>angle 0.0</gparam>
<lparam>ADDRESS_BITS 8</lparam>
<lparam>DATA_BITS 8</lparam></gate>
<gate>
<ID>33</ID>
<type>DD_KEYPAD_HEX</type>
<position>-10,40</position>
<output>
<ID>OUT_0</ID>113 </output>
<output>
<ID>OUT_1</ID>114 </output>
<output>
<ID>OUT_2</ID>115 </output>
<output>
<ID>OUT_3</ID>116 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 15</lparam></gate>
<gate>
<ID>34</ID>
<type>DD_KEYPAD_HEX</type>
<position>-22,40</position>
<output>
<ID>OUT_0</ID>117 </output>
<output>
<ID>OUT_1</ID>118 </output>
<output>
<ID>OUT_2</ID>119 </output>
<output>
<ID>OUT_3</ID>120 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 2</lparam></gate>
<gate>
<ID>35</ID>
<type>AA_TOGGLE</type>
<position>14.5,39.5</position>
<output>
<ID>OUT_0</ID>121 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>36</ID>
<type>AE_SMALL_INVERTER</type>
<position>-25.5,28</position>
<input>
<ID>IN_0</ID>9 </input>
<output>
<ID>OUT_0</ID>14 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>37</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>5,-5.5</position>
<input>
<ID>ENABLE_0</ID>121 </input>
<input>
<ID>IN_0</ID>15 </input>
<input>
<ID>IN_1</ID>16 </input>
<input>
<ID>IN_2</ID>17 </input>
<input>
<ID>IN_3</ID>18 </input>
<input>
<ID>IN_4</ID>26 </input>
<input>
<ID>IN_5</ID>27 </input>
<input>
<ID>IN_6</ID>28 </input>
<input>
<ID>IN_7</ID>37 </input>
<output>
<ID>OUT_0</ID>39 </output>
<output>
<ID>OUT_1</ID>38 </output>
<output>
<ID>OUT_2</ID>40 </output>
<output>
<ID>OUT_3</ID>41 </output>
<output>
<ID>OUT_4</ID>44 </output>
<output>
<ID>OUT_5</ID>45 </output>
<output>
<ID>OUT_6</ID>43 </output>
<output>
<ID>OUT_7</ID>42 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>38</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>5,-25.5</position>
<input>
<ID>ENABLE_0</ID>121 </input>
<input>
<ID>IN_0</ID>15 </input>
<input>
<ID>IN_1</ID>16 </input>
<input>
<ID>IN_2</ID>17 </input>
<input>
<ID>IN_3</ID>18 </input>
<input>
<ID>IN_4</ID>26 </input>
<input>
<ID>IN_5</ID>27 </input>
<input>
<ID>IN_6</ID>28 </input>
<input>
<ID>IN_7</ID>37 </input>
<output>
<ID>OUT_0</ID>53 </output>
<output>
<ID>OUT_1</ID>47 </output>
<output>
<ID>OUT_2</ID>46 </output>
<output>
<ID>OUT_3</ID>50 </output>
<output>
<ID>OUT_4</ID>48 </output>
<output>
<ID>OUT_5</ID>49 </output>
<output>
<ID>OUT_6</ID>51 </output>
<output>
<ID>OUT_7</ID>52 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>39</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>5,-46</position>
<input>
<ID>ENABLE_0</ID>121 </input>
<input>
<ID>IN_0</ID>15 </input>
<input>
<ID>IN_1</ID>16 </input>
<input>
<ID>IN_2</ID>17 </input>
<input>
<ID>IN_3</ID>18 </input>
<input>
<ID>IN_4</ID>26 </input>
<input>
<ID>IN_5</ID>27 </input>
<input>
<ID>IN_6</ID>28 </input>
<input>
<ID>IN_7</ID>37 </input>
<output>
<ID>OUT_0</ID>57 </output>
<output>
<ID>OUT_1</ID>61 </output>
<output>
<ID>OUT_2</ID>58 </output>
<output>
<ID>OUT_3</ID>54 </output>
<output>
<ID>OUT_4</ID>59 </output>
<output>
<ID>OUT_5</ID>55 </output>
<output>
<ID>OUT_6</ID>56 </output>
<output>
<ID>OUT_7</ID>60 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>40</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>5.5,-65</position>
<input>
<ID>ENABLE_0</ID>121 </input>
<input>
<ID>IN_0</ID>15 </input>
<input>
<ID>IN_1</ID>16 </input>
<input>
<ID>IN_2</ID>17 </input>
<input>
<ID>IN_3</ID>18 </input>
<input>
<ID>IN_4</ID>26 </input>
<input>
<ID>IN_5</ID>27 </input>
<input>
<ID>IN_6</ID>28 </input>
<input>
<ID>IN_7</ID>37 </input>
<output>
<ID>OUT_0</ID>64 </output>
<output>
<ID>OUT_1</ID>63 </output>
<output>
<ID>OUT_2</ID>69 </output>
<output>
<ID>OUT_3</ID>65 </output>
<output>
<ID>OUT_4</ID>66 </output>
<output>
<ID>OUT_5</ID>67 </output>
<output>
<ID>OUT_6</ID>62 </output>
<output>
<ID>OUT_7</ID>68 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>41</ID>
<type>AE_OR2</type>
<position>-3,15</position>
<input>
<ID>IN_0</ID>13 </input>
<input>
<ID>IN_1</ID>11 </input>
<output>
<ID>OUT</ID>70 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>42</ID>
<type>AE_FULLADDER_4BIT</type>
<position>81.5,-59</position>
<input>
<ID>IN_0</ID>81 </input>
<input>
<ID>IN_1</ID>82 </input>
<input>
<ID>IN_2</ID>83 </input>
<input>
<ID>IN_3</ID>84 </input>
<input>
<ID>IN_B_0</ID>77 </input>
<input>
<ID>IN_B_1</ID>78 </input>
<input>
<ID>IN_B_2</ID>79 </input>
<input>
<ID>IN_B_3</ID>80 </input>
<output>
<ID>OUT_0</ID>104 </output>
<output>
<ID>OUT_1</ID>105 </output>
<output>
<ID>OUT_2</ID>106 </output>
<output>
<ID>OUT_3</ID>107 </output>
<output>
<ID>carry_out</ID>76 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>43</ID>
<type>AE_FULLADDER_4BIT</type>
<position>96.5,-59.5</position>
<input>
<ID>IN_0</ID>89 </input>
<input>
<ID>IN_1</ID>90 </input>
<input>
<ID>IN_2</ID>91 </input>
<input>
<ID>IN_3</ID>92 </input>
<input>
<ID>IN_B_0</ID>85 </input>
<input>
<ID>IN_B_1</ID>86 </input>
<input>
<ID>IN_B_2</ID>87 </input>
<input>
<ID>IN_B_3</ID>88 </input>
<output>
<ID>OUT_0</ID>108 </output>
<output>
<ID>OUT_1</ID>109 </output>
<output>
<ID>OUT_2</ID>110 </output>
<output>
<ID>OUT_3</ID>111 </output>
<input>
<ID>carry_in</ID>76 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>44</ID>
<type>AA_AND2</type>
<position>83.5,-10</position>
<input>
<ID>IN_0</ID>88 </input>
<input>
<ID>IN_1</ID>92 </input>
<output>
<ID>OUT</ID>95 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>45</ID>
<type>AA_AND2</type>
<position>83.5,-14.5</position>
<input>
<ID>IN_0</ID>87 </input>
<input>
<ID>IN_1</ID>91 </input>
<output>
<ID>OUT</ID>96 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>46</ID>
<type>AA_AND2</type>
<position>83.5,-19</position>
<input>
<ID>IN_0</ID>86 </input>
<input>
<ID>IN_1</ID>90 </input>
<output>
<ID>OUT</ID>97 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>47</ID>
<type>AA_AND2</type>
<position>83.5,-23.5</position>
<input>
<ID>IN_0</ID>85 </input>
<input>
<ID>IN_1</ID>89 </input>
<output>
<ID>OUT</ID>98 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>48</ID>
<type>AA_AND2</type>
<position>83.5,-28</position>
<input>
<ID>IN_0</ID>80 </input>
<input>
<ID>IN_1</ID>84 </input>
<output>
<ID>OUT</ID>99 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>49</ID>
<type>AA_AND2</type>
<position>83.5,-32.5</position>
<input>
<ID>IN_0</ID>79 </input>
<input>
<ID>IN_1</ID>83 </input>
<output>
<ID>OUT</ID>100 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>50</ID>
<type>AA_AND2</type>
<position>83.5,-37</position>
<input>
<ID>IN_0</ID>78 </input>
<input>
<ID>IN_1</ID>82 </input>
<output>
<ID>OUT</ID>101 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>51</ID>
<type>AA_AND2</type>
<position>83.5,-41.5</position>
<input>
<ID>IN_0</ID>77 </input>
<input>
<ID>IN_1</ID>81 </input>
<output>
<ID>OUT</ID>102 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>52</ID>
<type>AA_MUX_2x1</type>
<position>102,-14.5</position>
<input>
<ID>IN_0</ID>111 </input>
<input>
<ID>IN_1</ID>95 </input>
<output>
<ID>OUT</ID>25 </output>
<input>
<ID>SEL_0</ID>112 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>53</ID>
<type>AA_MUX_2x1</type>
<position>102,-19</position>
<input>
<ID>IN_0</ID>110 </input>
<input>
<ID>IN_1</ID>96 </input>
<output>
<ID>OUT</ID>24 </output>
<input>
<ID>SEL_0</ID>112 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>54</ID>
<type>AA_MUX_2x1</type>
<position>102,-32.5</position>
<input>
<ID>IN_0</ID>107 </input>
<input>
<ID>IN_1</ID>99 </input>
<output>
<ID>OUT</ID>21 </output>
<input>
<ID>SEL_0</ID>112 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>55</ID>
<type>AA_MUX_2x1</type>
<position>102,-37</position>
<input>
<ID>IN_0</ID>106 </input>
<input>
<ID>IN_1</ID>100 </input>
<output>
<ID>OUT</ID>20 </output>
<input>
<ID>SEL_0</ID>112 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>56</ID>
<type>AA_MUX_2x1</type>
<position>102,-28</position>
<input>
<ID>IN_0</ID>108 </input>
<input>
<ID>IN_1</ID>98 </input>
<output>
<ID>OUT</ID>22 </output>
<input>
<ID>SEL_0</ID>112 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>57</ID>
<type>AA_MUX_2x1</type>
<position>102,-23.5</position>
<input>
<ID>IN_0</ID>109 </input>
<input>
<ID>IN_1</ID>97 </input>
<output>
<ID>OUT</ID>23 </output>
<input>
<ID>SEL_0</ID>112 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>58</ID>
<type>AA_MUX_2x1</type>
<position>102,-46</position>
<input>
<ID>IN_0</ID>104 </input>
<input>
<ID>IN_1</ID>102 </input>
<output>
<ID>OUT</ID>103 </output>
<input>
<ID>SEL_0</ID>112 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>59</ID>
<type>AA_MUX_2x1</type>
<position>102,-41.5</position>
<input>
<ID>IN_0</ID>105 </input>
<input>
<ID>IN_1</ID>101 </input>
<output>
<ID>OUT</ID>19 </output>
<input>
<ID>SEL_0</ID>112 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>60</ID>
<type>AE_REGISTER8</type>
<position>15,-6</position>
<input>
<ID>IN_0</ID>39 </input>
<input>
<ID>IN_1</ID>38 </input>
<input>
<ID>IN_2</ID>40 </input>
<input>
<ID>IN_3</ID>41 </input>
<input>
<ID>IN_4</ID>44 </input>
<input>
<ID>IN_5</ID>45 </input>
<input>
<ID>IN_6</ID>43 </input>
<input>
<ID>IN_7</ID>42 </input>
<output>
<ID>OUT_0</ID>133 </output>
<output>
<ID>OUT_1</ID>133 </output>
<output>
<ID>OUT_2</ID>131 </output>
<output>
<ID>OUT_3</ID>130 </output>
<output>
<ID>OUT_4</ID>129 </output>
<output>
<ID>OUT_5</ID>128 </output>
<output>
<ID>OUT_6</ID>127 </output>
<output>
<ID>OUT_7</ID>126 </output>
<input>
<ID>clock</ID>75 </input>
<input>
<ID>load</ID>74 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 9</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>61</ID>
<type>BB_CLOCK</type>
<position>-27.5,-78.5</position>
<output>
<ID>CLK</ID>75 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>62</ID>
<type>AE_MUX_4x1</type>
<position>38,-1</position>
<input>
<ID>IN_0</ID>8 </input>
<input>
<ID>IN_1</ID>142 </input>
<input>
<ID>IN_2</ID>134 </input>
<input>
<ID>IN_3</ID>126 </input>
<output>
<ID>OUT</ID>88 </output>
<input>
<ID>SEL_0</ID>94 </input>
<input>
<ID>SEL_1</ID>93 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<wire>
<ID>1</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>19,-76.5,45,-76.5</points>
<connection>
<GID>14</GID>
<name>IN_0</name></connection>
<connection>
<GID>7</GID>
<name>IN_0</name></connection>
<intersection>19 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>19,-76.5,19,-68.5</points>
<connection>
<GID>24</GID>
<name>OUT_0</name></connection>
<intersection>-76.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>19,-67.5,45,-67.5</points>
<connection>
<GID>24</GID>
<name>OUT_1</name></connection>
<intersection>35 13</intersection>
<intersection>45 14</intersection></hsegment>
<vsegment>
<ID>13</ID>
<points>35,-67.5,35,-66.5</points>
<connection>
<GID>6</GID>
<name>IN_0</name></connection>
<intersection>-67.5 1</intersection></vsegment>
<vsegment>
<ID>14</ID>
<points>45,-67.5,45,-66.5</points>
<connection>
<GID>13</GID>
<name>IN_0</name></connection>
<intersection>-67.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>29,-56.5,45,-56.5</points>
<connection>
<GID>12</GID>
<name>IN_0</name></connection>
<connection>
<GID>5</GID>
<name>IN_0</name></connection>
<intersection>29 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>29,-66.5,29,-56.5</points>
<intersection>-66.5 4</intersection>
<intersection>-56.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>19,-66.5,29,-66.5</points>
<connection>
<GID>24</GID>
<name>OUT_2</name></connection>
<intersection>29 3</intersection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>28,-46,45,-46</points>
<connection>
<GID>11</GID>
<name>IN_0</name></connection>
<intersection>28 3</intersection>
<intersection>35 15</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>28,-65.5,28,-46</points>
<intersection>-65.5 4</intersection>
<intersection>-46 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>19,-65.5,28,-65.5</points>
<connection>
<GID>24</GID>
<name>OUT_3</name></connection>
<intersection>28 3</intersection></hsegment>
<vsegment>
<ID>15</ID>
<points>35,-46.5,35,-46</points>
<connection>
<GID>4</GID>
<name>IN_0</name></connection>
<intersection>-46 1</intersection></vsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>27,-36,45,-36</points>
<connection>
<GID>10</GID>
<name>IN_0</name></connection>
<connection>
<GID>3</GID>
<name>IN_0</name></connection>
<intersection>27 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>27,-64.5,27,-36</points>
<intersection>-64.5 4</intersection>
<intersection>-36 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>19,-64.5,27,-64.5</points>
<connection>
<GID>24</GID>
<name>OUT_4</name></connection>
<intersection>27 3</intersection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>26,-25,45,-25</points>
<connection>
<GID>9</GID>
<name>IN_0</name></connection>
<connection>
<GID>2</GID>
<name>IN_0</name></connection>
<intersection>26 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>26,-63.5,26,-25</points>
<intersection>-63.5 4</intersection>
<intersection>-25 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>19,-63.5,26,-63.5</points>
<connection>
<GID>24</GID>
<name>OUT_5</name></connection>
<intersection>26 3</intersection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>24.5,-14,45,-14</points>
<connection>
<GID>8</GID>
<name>IN_0</name></connection>
<connection>
<GID>1</GID>
<name>IN_0</name></connection>
<intersection>24.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>24.5,-62.5,24.5,-14</points>
<intersection>-62.5 4</intersection>
<intersection>-14 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>19,-62.5,24.5,-62.5</points>
<connection>
<GID>24</GID>
<name>OUT_6</name></connection>
<intersection>24.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>23,-4,45,-4</points>
<connection>
<GID>62</GID>
<name>IN_0</name></connection>
<connection>
<GID>15</GID>
<name>IN_0</name></connection>
<intersection>23 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>23,-61.5,23,-4</points>
<intersection>-61.5 4</intersection>
<intersection>-4 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>19,-61.5,23,-61.5</points>
<connection>
<GID>24</GID>
<name>OUT_7</name></connection>
<intersection>23 3</intersection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-27.5,17.5,21,17.5</points>
<intersection>-27.5 6</intersection>
<intersection>-8.5 3</intersection>
<intersection>21 7</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-8.5,17.5,-8.5,19.5</points>
<intersection>17.5 1</intersection>
<intersection>19.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-12.5,19.5,-8.5,19.5</points>
<connection>
<GID>27</GID>
<name>OUT_0</name></connection>
<intersection>-8.5 3</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>-27.5,14.5,-27.5,28</points>
<connection>
<GID>36</GID>
<name>IN_0</name></connection>
<intersection>14.5 12</intersection>
<intersection>17.5 1</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>21,10,21,17.5</points>
<intersection>10 9</intersection>
<intersection>17.5 1</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>21,10,61.5,10</points>
<intersection>21 7</intersection>
<intersection>55.5 14</intersection>
<intersection>61.5 13</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>-30.5,14.5,-27.5,14.5</points>
<connection>
<GID>31</GID>
<name>write_enable</name></connection>
<intersection>-27.5 6</intersection></hsegment>
<vsegment>
<ID>13</ID>
<points>61.5,9.5,61.5,10</points>
<connection>
<GID>16</GID>
<name>ENABLE_0</name></connection>
<intersection>10 9</intersection></vsegment>
<vsegment>
<ID>14</ID>
<points>55.5,10,55.5,26.5</points>
<intersection>10 9</intersection>
<intersection>23.5 18</intersection>
<intersection>26.5 22</intersection></vsegment>
<hsegment>
<ID>18</ID>
<points>44.5,23.5,55.5,23.5</points>
<intersection>44.5 20</intersection>
<intersection>55.5 14</intersection></hsegment>
<vsegment>
<ID>20</ID>
<points>44.5,23.5,44.5,26.5</points>
<connection>
<GID>20</GID>
<name>ENABLE_0</name></connection>
<intersection>23.5 18</intersection></vsegment>
<hsegment>
<ID>22</ID>
<points>55,26.5,55.5,26.5</points>
<connection>
<GID>18</GID>
<name>IN_0</name></connection>
<intersection>55.5 14</intersection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-7.5,13.5,-7.5,20.5</points>
<intersection>13.5 1</intersection>
<intersection>20.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-30.5,13.5,-7.5,13.5</points>
<connection>
<GID>31</GID>
<name>ENABLE_0</name></connection>
<intersection>-26 3</intersection>
<intersection>-7.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-12.5,20.5,-7.5,20.5</points>
<connection>
<GID>27</GID>
<name>OUT_1</name></connection>
<intersection>-7.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-26,-20.5,-26,13.5</points>
<connection>
<GID>21</GID>
<name>ENABLE_0</name></connection>
<intersection>13.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>101,-1,101,21.5</points>
<connection>
<GID>29</GID>
<name>IN_0</name></connection>
<intersection>21.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-12.5,21.5,101,21.5</points>
<connection>
<GID>27</GID>
<name>OUT_2</name></connection>
<intersection>-3 2</intersection>
<intersection>101 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-3,18,-3,21.5</points>
<intersection>18 6</intersection>
<intersection>21.5 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>-4,18,-3,18</points>
<connection>
<GID>41</GID>
<name>IN_1</name></connection>
<intersection>-3 2</intersection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<vsegment>
<ID>4</ID>
<points>101,-5.5,101,-5</points>
<connection>
<GID>30</GID>
<name>IN_1</name></connection>
<connection>
<GID>29</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>103,-5.5,103,22.5</points>
<connection>
<GID>30</GID>
<name>IN_0</name></connection>
<intersection>22.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-12.5,22.5,103,22.5</points>
<connection>
<GID>27</GID>
<name>OUT_3</name></connection>
<intersection>-2 3</intersection>
<intersection>103 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-2,18,-2,22.5</points>
<connection>
<GID>41</GID>
<name>IN_0</name></connection>
<intersection>22.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-23.5,28,-18.5,28</points>
<connection>
<GID>36</GID>
<name>OUT_0</name></connection>
<connection>
<GID>25</GID>
<name>ENABLE</name></connection></hsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-15.5,-68.5,-15.5,-9</points>
<intersection>-68.5 11</intersection>
<intersection>-49.5 9</intersection>
<intersection>-40.5 2</intersection>
<intersection>-29 6</intersection>
<intersection>-9 7</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-24,-40.5,-15.5,-40.5</points>
<connection>
<GID>19</GID>
<name>OUT_0</name></connection>
<intersection>-15.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-24,-29,3,-29</points>
<connection>
<GID>38</GID>
<name>IN_0</name></connection>
<connection>
<GID>21</GID>
<name>OUT_0</name></connection>
<intersection>-15.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-15.5,-9,3,-9</points>
<connection>
<GID>37</GID>
<name>IN_0</name></connection>
<intersection>-15.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>-15.5,-49.5,3,-49.5</points>
<connection>
<GID>39</GID>
<name>IN_0</name></connection>
<intersection>-15.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>-15.5,-68.5,3.5,-68.5</points>
<connection>
<GID>40</GID>
<name>IN_0</name></connection>
<intersection>-15.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-14.5,-67.5,-14.5,-8</points>
<intersection>-67.5 16</intersection>
<intersection>-48.5 14</intersection>
<intersection>-39.5 2</intersection>
<intersection>-28 5</intersection>
<intersection>-8 13</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-24,-39.5,-14.5,-39.5</points>
<connection>
<GID>19</GID>
<name>OUT_1</name></connection>
<intersection>-14.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-24,-28,3,-28</points>
<connection>
<GID>38</GID>
<name>IN_1</name></connection>
<connection>
<GID>21</GID>
<name>OUT_1</name></connection>
<intersection>-14.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>-14.5,-8,3,-8</points>
<connection>
<GID>37</GID>
<name>IN_1</name></connection>
<intersection>-14.5 0</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>-14.5,-48.5,3,-48.5</points>
<connection>
<GID>39</GID>
<name>IN_1</name></connection>
<intersection>-14.5 0</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>-14.5,-67.5,3.5,-67.5</points>
<connection>
<GID>40</GID>
<name>IN_1</name></connection>
<intersection>-14.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-13.5,-66.5,-13.5,-7</points>
<intersection>-66.5 15</intersection>
<intersection>-47.5 13</intersection>
<intersection>-38.5 2</intersection>
<intersection>-27 4</intersection>
<intersection>-7 12</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-24,-38.5,-13.5,-38.5</points>
<connection>
<GID>19</GID>
<name>OUT_2</name></connection>
<intersection>-13.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-24,-27,3,-27</points>
<connection>
<GID>38</GID>
<name>IN_2</name></connection>
<connection>
<GID>21</GID>
<name>OUT_2</name></connection>
<intersection>-13.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>-13.5,-7,3,-7</points>
<connection>
<GID>37</GID>
<name>IN_2</name></connection>
<intersection>-13.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>-13.5,-47.5,3,-47.5</points>
<connection>
<GID>39</GID>
<name>IN_2</name></connection>
<intersection>-13.5 0</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>-13.5,-66.5,3.5,-66.5</points>
<connection>
<GID>40</GID>
<name>IN_2</name></connection>
<intersection>-13.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-12.5,-65.5,-12.5,-6</points>
<intersection>-65.5 9</intersection>
<intersection>-46.5 7</intersection>
<intersection>-37.5 2</intersection>
<intersection>-26 4</intersection>
<intersection>-6 6</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-24,-37.5,-12.5,-37.5</points>
<connection>
<GID>19</GID>
<name>OUT_3</name></connection>
<intersection>-12.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-24,-26,3,-26</points>
<connection>
<GID>38</GID>
<name>IN_3</name></connection>
<connection>
<GID>21</GID>
<name>OUT_3</name></connection>
<intersection>-12.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-12.5,-6,3,-6</points>
<connection>
<GID>37</GID>
<name>IN_3</name></connection>
<intersection>-12.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-12.5,-46.5,3,-46.5</points>
<connection>
<GID>39</GID>
<name>IN_3</name></connection>
<intersection>-12.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>-12.5,-65.5,3.5,-65.5</points>
<connection>
<GID>40</GID>
<name>IN_3</name></connection>
<intersection>-12.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>105.5,-83,105.5,-41.5</points>
<intersection>-83 1</intersection>
<intersection>-41.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-34,-83,105.5,-83</points>
<intersection>-34 3</intersection>
<intersection>105.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>104,-41.5,105.5,-41.5</points>
<connection>
<GID>59</GID>
<name>OUT</name></connection>
<intersection>105.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-34,-83,-34,-39.5</points>
<intersection>-83 1</intersection>
<intersection>-39.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-34,-39.5,-28,-39.5</points>
<connection>
<GID>19</GID>
<name>IN_1</name></connection>
<intersection>-34 3</intersection></hsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>106.5,-84,106.5,-37</points>
<intersection>-84 1</intersection>
<intersection>-37 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-35,-84,106.5,-84</points>
<intersection>-35 3</intersection>
<intersection>106.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>104,-37,106.5,-37</points>
<connection>
<GID>55</GID>
<name>OUT</name></connection>
<intersection>106.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-35,-84,-35,-38.5</points>
<intersection>-84 1</intersection>
<intersection>-38.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>-35,-38.5,-28,-38.5</points>
<connection>
<GID>19</GID>
<name>IN_2</name></connection>
<intersection>-35 3</intersection></hsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>107.5,-85,107.5,-32.5</points>
<intersection>-85 1</intersection>
<intersection>-32.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-36,-85,107.5,-85</points>
<intersection>-36 3</intersection>
<intersection>107.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>104,-32.5,107.5,-32.5</points>
<connection>
<GID>54</GID>
<name>OUT</name></connection>
<intersection>107.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-36,-85,-36,-37.5</points>
<intersection>-85 1</intersection>
<intersection>-37.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-36,-37.5,-28,-37.5</points>
<connection>
<GID>19</GID>
<name>IN_3</name></connection>
<intersection>-36 3</intersection></hsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>108.5,-86,108.5,-28</points>
<intersection>-86 1</intersection>
<intersection>-28 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-37,-86,108.5,-86</points>
<intersection>-37 3</intersection>
<intersection>108.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>104,-28,108.5,-28</points>
<connection>
<GID>56</GID>
<name>OUT</name></connection>
<intersection>108.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-37,-86,-37,-36.5</points>
<intersection>-86 1</intersection>
<intersection>-36.5 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>-37,-36.5,-28,-36.5</points>
<connection>
<GID>19</GID>
<name>IN_4</name></connection>
<intersection>-37 3</intersection></hsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>109.5,-87,109.5,-23.5</points>
<intersection>-87 1</intersection>
<intersection>-23.5 9</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-38,-87,109.5,-87</points>
<intersection>-38 3</intersection>
<intersection>109.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-38,-87,-38,-35.5</points>
<intersection>-87 1</intersection>
<intersection>-35.5 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>-38,-35.5,-28,-35.5</points>
<connection>
<GID>19</GID>
<name>IN_5</name></connection>
<intersection>-38 3</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>104,-23.5,109.5,-23.5</points>
<connection>
<GID>57</GID>
<name>OUT</name></connection>
<intersection>109.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>24</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>110.5,-88,110.5,-19</points>
<intersection>-88 1</intersection>
<intersection>-19 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-39,-88,110.5,-88</points>
<intersection>-39 3</intersection>
<intersection>110.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>104,-19,110.5,-19</points>
<connection>
<GID>53</GID>
<name>OUT</name></connection>
<intersection>110.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-39,-88,-39,-34.5</points>
<intersection>-88 1</intersection>
<intersection>-34.5 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>-39,-34.5,-28,-34.5</points>
<connection>
<GID>19</GID>
<name>IN_6</name></connection>
<intersection>-39 3</intersection></hsegment></shape></wire>
<wire>
<ID>25</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>111.5,-89,111.5,-14.5</points>
<intersection>-89 1</intersection>
<intersection>-14.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-40,-89,111.5,-89</points>
<intersection>-40 3</intersection>
<intersection>111.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>104,-14.5,111.5,-14.5</points>
<connection>
<GID>52</GID>
<name>OUT</name></connection>
<intersection>111.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-40,-89,-40,-33.5</points>
<intersection>-89 1</intersection>
<intersection>-33.5 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>-40,-33.5,-28,-33.5</points>
<connection>
<GID>19</GID>
<name>IN_7</name></connection>
<intersection>-40 3</intersection></hsegment></shape></wire>
<wire>
<ID>26</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-11.5,-64.5,-11.5,-5</points>
<intersection>-64.5 14</intersection>
<intersection>-45.5 12</intersection>
<intersection>-36.5 2</intersection>
<intersection>-25 4</intersection>
<intersection>-5 11</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-24,-36.5,-11.5,-36.5</points>
<connection>
<GID>19</GID>
<name>OUT_4</name></connection>
<intersection>-11.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-24,-25,3,-25</points>
<connection>
<GID>38</GID>
<name>IN_4</name></connection>
<connection>
<GID>21</GID>
<name>OUT_4</name></connection>
<intersection>-11.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>-11.5,-5,3,-5</points>
<connection>
<GID>37</GID>
<name>IN_4</name></connection>
<intersection>-11.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>-11.5,-45.5,3,-45.5</points>
<connection>
<GID>39</GID>
<name>IN_4</name></connection>
<intersection>-11.5 0</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>-11.5,-64.5,3.5,-64.5</points>
<connection>
<GID>40</GID>
<name>IN_4</name></connection>
<intersection>-11.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>27</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-10.5,-63.5,-10.5,-4</points>
<intersection>-63.5 14</intersection>
<intersection>-44.5 12</intersection>
<intersection>-35.5 2</intersection>
<intersection>-24 4</intersection>
<intersection>-4 11</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-24,-35.5,-10.5,-35.5</points>
<connection>
<GID>19</GID>
<name>OUT_5</name></connection>
<intersection>-10.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-24,-24,3,-24</points>
<connection>
<GID>38</GID>
<name>IN_5</name></connection>
<connection>
<GID>21</GID>
<name>OUT_5</name></connection>
<intersection>-10.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>-10.5,-4,3,-4</points>
<connection>
<GID>37</GID>
<name>IN_5</name></connection>
<intersection>-10.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>-10.5,-44.5,3,-44.5</points>
<connection>
<GID>39</GID>
<name>IN_5</name></connection>
<intersection>-10.5 0</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>-10.5,-63.5,3.5,-63.5</points>
<connection>
<GID>40</GID>
<name>IN_5</name></connection>
<intersection>-10.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>28</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-9.5,-62.5,-9.5,-3</points>
<intersection>-62.5 18</intersection>
<intersection>-43.5 16</intersection>
<intersection>-34.5 2</intersection>
<intersection>-23 4</intersection>
<intersection>-3 15</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-24,-34.5,-9.5,-34.5</points>
<connection>
<GID>19</GID>
<name>OUT_6</name></connection>
<intersection>-9.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-24,-23,3,-23</points>
<connection>
<GID>38</GID>
<name>IN_6</name></connection>
<connection>
<GID>21</GID>
<name>OUT_6</name></connection>
<intersection>-9.5 0</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>-9.5,-3,3,-3</points>
<connection>
<GID>37</GID>
<name>IN_6</name></connection>
<intersection>-9.5 0</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>-9.5,-43.5,3,-43.5</points>
<connection>
<GID>39</GID>
<name>IN_6</name></connection>
<intersection>-9.5 0</intersection></hsegment>
<hsegment>
<ID>18</ID>
<points>-9.5,-62.5,3.5,-62.5</points>
<connection>
<GID>40</GID>
<name>IN_6</name></connection>
<intersection>-9.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>29</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-32,-29,-32,7</points>
<connection>
<GID>31</GID>
<name>DATA_OUT_0</name></connection>
<connection>
<GID>31</GID>
<name>DATA_IN_0</name></connection>
<intersection>-29 5</intersection>
<intersection>1.5 6</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-32,-29,-28,-29</points>
<connection>
<GID>21</GID>
<name>IN_0</name></connection>
<intersection>-32 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-32,1.5,14,1.5</points>
<intersection>-32 0</intersection>
<intersection>14 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>14,1.5,14,12</points>
<intersection>1.5 6</intersection>
<intersection>12 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>14,12,67,12</points>
<intersection>14 7</intersection>
<intersection>67 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>67,1,67,12</points>
<intersection>1 10</intersection>
<intersection>12 8</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>63.5,1,67,1</points>
<connection>
<GID>16</GID>
<name>OUT_0</name></connection>
<intersection>67 9</intersection></hsegment></shape></wire>
<wire>
<ID>30</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-33,-28,-33,7</points>
<connection>
<GID>31</GID>
<name>DATA_OUT_1</name></connection>
<connection>
<GID>31</GID>
<name>DATA_IN_1</name></connection>
<intersection>-28 13</intersection>
<intersection>2 14</intersection></vsegment>
<hsegment>
<ID>13</ID>
<points>-33,-28,-28,-28</points>
<connection>
<GID>21</GID>
<name>IN_1</name></connection>
<intersection>-33 0</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>-33,2,13.5,2</points>
<intersection>-33 0</intersection>
<intersection>13.5 15</intersection></hsegment>
<vsegment>
<ID>15</ID>
<points>13.5,2,13.5,12.5</points>
<intersection>2 14</intersection>
<intersection>12.5 16</intersection></vsegment>
<hsegment>
<ID>16</ID>
<points>13.5,12.5,66.5,12.5</points>
<intersection>13.5 15</intersection>
<intersection>66.5 17</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>66.5,2,66.5,12.5</points>
<intersection>2 18</intersection>
<intersection>12.5 16</intersection></vsegment>
<hsegment>
<ID>18</ID>
<points>63.5,2,66.5,2</points>
<connection>
<GID>16</GID>
<name>OUT_1</name></connection>
<intersection>66.5 17</intersection></hsegment></shape></wire>
<wire>
<ID>31</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-34,-27,-34,7</points>
<connection>
<GID>31</GID>
<name>DATA_OUT_2</name></connection>
<connection>
<GID>31</GID>
<name>DATA_IN_2</name></connection>
<intersection>-27 1</intersection>
<intersection>2.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-34,-27,-28,-27</points>
<connection>
<GID>21</GID>
<name>IN_2</name></connection>
<intersection>-34 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-34,2.5,13,2.5</points>
<intersection>-34 0</intersection>
<intersection>13 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>13,2.5,13,13</points>
<intersection>2.5 3</intersection>
<intersection>13 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>13,13,66,13</points>
<intersection>13 4</intersection>
<intersection>66 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>66,3,66,13</points>
<intersection>3 7</intersection>
<intersection>13 5</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>63.5,3,66,3</points>
<connection>
<GID>16</GID>
<name>OUT_2</name></connection>
<intersection>66 6</intersection></hsegment></shape></wire>
<wire>
<ID>32</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-35,-26,-35,7</points>
<connection>
<GID>31</GID>
<name>DATA_OUT_3</name></connection>
<connection>
<GID>31</GID>
<name>DATA_IN_3</name></connection>
<intersection>-26 1</intersection>
<intersection>3 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-35,-26,-28,-26</points>
<connection>
<GID>21</GID>
<name>IN_3</name></connection>
<intersection>-35 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-35,3,12.5,3</points>
<intersection>-35 0</intersection>
<intersection>12.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>12.5,3,12.5,13.5</points>
<intersection>3 3</intersection>
<intersection>13.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>12.5,13.5,65.5,13.5</points>
<intersection>12.5 4</intersection>
<intersection>65.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>65.5,4,65.5,13.5</points>
<intersection>4 7</intersection>
<intersection>13.5 5</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>63.5,4,65.5,4</points>
<connection>
<GID>16</GID>
<name>OUT_3</name></connection>
<intersection>65.5 6</intersection></hsegment></shape></wire>
<wire>
<ID>33</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-36,-25,-36,7</points>
<connection>
<GID>31</GID>
<name>DATA_OUT_4</name></connection>
<connection>
<GID>31</GID>
<name>DATA_IN_4</name></connection>
<intersection>-25 1</intersection>
<intersection>3.5 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-36,-25,-28,-25</points>
<connection>
<GID>21</GID>
<name>IN_4</name></connection>
<intersection>-36 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-36,3.5,12,3.5</points>
<intersection>-36 0</intersection>
<intersection>12 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>12,3.5,12,14</points>
<intersection>3.5 4</intersection>
<intersection>14 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>12,14,65,14</points>
<intersection>12 5</intersection>
<intersection>65 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>65,5,65,14</points>
<intersection>5 8</intersection>
<intersection>14 6</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>63.5,5,65,5</points>
<connection>
<GID>16</GID>
<name>OUT_4</name></connection>
<intersection>65 7</intersection></hsegment></shape></wire>
<wire>
<ID>34</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-37,-24,-37,7</points>
<connection>
<GID>31</GID>
<name>DATA_OUT_5</name></connection>
<connection>
<GID>31</GID>
<name>DATA_IN_5</name></connection>
<intersection>-24 1</intersection>
<intersection>4 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-37,-24,-28,-24</points>
<connection>
<GID>21</GID>
<name>IN_5</name></connection>
<intersection>-37 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-37,4,11.5,4</points>
<intersection>-37 0</intersection>
<intersection>11.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>11.5,4,11.5,14.5</points>
<intersection>4 3</intersection>
<intersection>14.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>11.5,14.5,64.5,14.5</points>
<intersection>11.5 4</intersection>
<intersection>64.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>64.5,6,64.5,14.5</points>
<intersection>6 7</intersection>
<intersection>14.5 5</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>63.5,6,64.5,6</points>
<connection>
<GID>16</GID>
<name>OUT_5</name></connection>
<intersection>64.5 6</intersection></hsegment></shape></wire>
<wire>
<ID>35</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-38,-23,-38,7</points>
<connection>
<GID>31</GID>
<name>DATA_OUT_6</name></connection>
<connection>
<GID>31</GID>
<name>DATA_IN_6</name></connection>
<intersection>-23 1</intersection>
<intersection>4.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-38,-23,-28,-23</points>
<connection>
<GID>21</GID>
<name>IN_6</name></connection>
<intersection>-38 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-38,4.5,11,4.5</points>
<intersection>-38 0</intersection>
<intersection>11 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>11,4.5,11,15</points>
<intersection>4.5 3</intersection>
<intersection>15 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>11,15,64,15</points>
<intersection>11 4</intersection>
<intersection>64 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>64,7,64,15</points>
<intersection>7 7</intersection>
<intersection>15 5</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>63.5,7,64,7</points>
<connection>
<GID>16</GID>
<name>OUT_6</name></connection>
<intersection>64 6</intersection></hsegment></shape></wire>
<wire>
<ID>36</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-39,-22,-39,7</points>
<connection>
<GID>31</GID>
<name>DATA_OUT_7</name></connection>
<connection>
<GID>31</GID>
<name>DATA_IN_7</name></connection>
<intersection>-22 1</intersection>
<intersection>5 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-39,-22,-28,-22</points>
<connection>
<GID>21</GID>
<name>IN_7</name></connection>
<intersection>-39 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-39,5,10.5,5</points>
<intersection>-39 0</intersection>
<intersection>10.5 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>10.5,5,10.5,15.5</points>
<intersection>5 4</intersection>
<intersection>15.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>10.5,15.5,63.5,15.5</points>
<intersection>10.5 5</intersection>
<intersection>63.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>63.5,8,63.5,15.5</points>
<connection>
<GID>16</GID>
<name>OUT_7</name></connection>
<intersection>15.5 6</intersection></vsegment></shape></wire>
<wire>
<ID>37</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-8.5,-61.5,-8.5,-2</points>
<intersection>-61.5 8</intersection>
<intersection>-42.5 6</intersection>
<intersection>-33.5 4</intersection>
<intersection>-22 1</intersection>
<intersection>-2 5</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-24,-22,3,-22</points>
<connection>
<GID>38</GID>
<name>IN_7</name></connection>
<connection>
<GID>21</GID>
<name>OUT_7</name></connection>
<intersection>-8.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-24,-33.5,-8.5,-33.5</points>
<connection>
<GID>19</GID>
<name>OUT_7</name></connection>
<intersection>-8.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-8.5,-2,3,-2</points>
<connection>
<GID>37</GID>
<name>IN_7</name></connection>
<intersection>-8.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-8.5,-42.5,3,-42.5</points>
<connection>
<GID>39</GID>
<name>IN_7</name></connection>
<intersection>-8.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-8.5,-61.5,3.5,-61.5</points>
<connection>
<GID>40</GID>
<name>IN_7</name></connection>
<intersection>-8.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>38</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>7,-8,11,-8</points>
<connection>
<GID>60</GID>
<name>IN_1</name></connection>
<connection>
<GID>37</GID>
<name>OUT_1</name></connection></hsegment></shape></wire>
<wire>
<ID>39</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>7,-9,11,-9</points>
<connection>
<GID>60</GID>
<name>IN_0</name></connection>
<connection>
<GID>37</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>40</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>7,-7,11,-7</points>
<connection>
<GID>60</GID>
<name>IN_2</name></connection>
<connection>
<GID>37</GID>
<name>OUT_2</name></connection></hsegment></shape></wire>
<wire>
<ID>41</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>7,-6,11,-6</points>
<connection>
<GID>60</GID>
<name>IN_3</name></connection>
<connection>
<GID>37</GID>
<name>OUT_3</name></connection></hsegment></shape></wire>
<wire>
<ID>42</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>7,-2,11,-2</points>
<connection>
<GID>60</GID>
<name>IN_7</name></connection>
<connection>
<GID>37</GID>
<name>OUT_7</name></connection></hsegment></shape></wire>
<wire>
<ID>43</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>7,-3,11,-3</points>
<connection>
<GID>60</GID>
<name>IN_6</name></connection>
<connection>
<GID>37</GID>
<name>OUT_6</name></connection></hsegment></shape></wire>
<wire>
<ID>44</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>7,-5,11,-5</points>
<connection>
<GID>60</GID>
<name>IN_4</name></connection>
<connection>
<GID>37</GID>
<name>OUT_4</name></connection></hsegment></shape></wire>
<wire>
<ID>45</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>7,-4,11,-4</points>
<connection>
<GID>60</GID>
<name>IN_5</name></connection>
<connection>
<GID>37</GID>
<name>OUT_5</name></connection></hsegment></shape></wire>
<wire>
<ID>46</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>7,-27,11,-27</points>
<connection>
<GID>38</GID>
<name>OUT_2</name></connection>
<connection>
<GID>22</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>47</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>7,-28,11,-28</points>
<connection>
<GID>38</GID>
<name>OUT_1</name></connection>
<connection>
<GID>22</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>48</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>7,-25,11,-25</points>
<connection>
<GID>38</GID>
<name>OUT_4</name></connection>
<connection>
<GID>22</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>49</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>7,-24,11,-24</points>
<connection>
<GID>38</GID>
<name>OUT_5</name></connection>
<connection>
<GID>22</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>50</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>7,-26,11,-26</points>
<connection>
<GID>38</GID>
<name>OUT_3</name></connection>
<connection>
<GID>22</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>51</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>7,-23,11,-23</points>
<connection>
<GID>38</GID>
<name>OUT_6</name></connection>
<connection>
<GID>22</GID>
<name>IN_6</name></connection></hsegment></shape></wire>
<wire>
<ID>52</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>7,-22,11,-22</points>
<connection>
<GID>38</GID>
<name>OUT_7</name></connection>
<connection>
<GID>22</GID>
<name>IN_7</name></connection></hsegment></shape></wire>
<wire>
<ID>53</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>7,-29,11,-29</points>
<connection>
<GID>38</GID>
<name>OUT_0</name></connection>
<connection>
<GID>22</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>54</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>7,-46.5,11,-46.5</points>
<connection>
<GID>39</GID>
<name>OUT_3</name></connection>
<connection>
<GID>23</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>55</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>7,-44.5,11,-44.5</points>
<connection>
<GID>39</GID>
<name>OUT_5</name></connection>
<connection>
<GID>23</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>56</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>7,-43.5,11,-43.5</points>
<connection>
<GID>39</GID>
<name>OUT_6</name></connection>
<connection>
<GID>23</GID>
<name>IN_6</name></connection></hsegment></shape></wire>
<wire>
<ID>57</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>7,-49.5,11,-49.5</points>
<connection>
<GID>39</GID>
<name>OUT_0</name></connection>
<connection>
<GID>23</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>58</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>7,-47.5,11,-47.5</points>
<connection>
<GID>39</GID>
<name>OUT_2</name></connection>
<connection>
<GID>23</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>59</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>7,-45.5,11,-45.5</points>
<connection>
<GID>39</GID>
<name>OUT_4</name></connection>
<connection>
<GID>23</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>60</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>7,-42.5,11,-42.5</points>
<connection>
<GID>39</GID>
<name>OUT_7</name></connection>
<connection>
<GID>23</GID>
<name>IN_7</name></connection></hsegment></shape></wire>
<wire>
<ID>61</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>7,-48.5,11,-48.5</points>
<connection>
<GID>39</GID>
<name>OUT_1</name></connection>
<connection>
<GID>23</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>62</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>7.5,-62.5,11,-62.5</points>
<connection>
<GID>40</GID>
<name>OUT_6</name></connection>
<connection>
<GID>24</GID>
<name>IN_6</name></connection></hsegment></shape></wire>
<wire>
<ID>63</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>7.5,-67.5,11,-67.5</points>
<connection>
<GID>40</GID>
<name>OUT_1</name></connection>
<connection>
<GID>24</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>64</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>7.5,-68.5,11,-68.5</points>
<connection>
<GID>40</GID>
<name>OUT_0</name></connection>
<connection>
<GID>24</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>65</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>7.5,-65.5,11,-65.5</points>
<connection>
<GID>40</GID>
<name>OUT_3</name></connection>
<connection>
<GID>24</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>66</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>7.5,-64.5,11,-64.5</points>
<connection>
<GID>40</GID>
<name>OUT_4</name></connection>
<connection>
<GID>24</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>67</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>7.5,-63.5,11,-63.5</points>
<connection>
<GID>40</GID>
<name>OUT_5</name></connection>
<connection>
<GID>24</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>68</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>7.5,-61.5,11,-61.5</points>
<connection>
<GID>40</GID>
<name>OUT_7</name></connection>
<connection>
<GID>24</GID>
<name>IN_7</name></connection></hsegment></shape></wire>
<wire>
<ID>69</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>7.5,-66.5,11,-66.5</points>
<connection>
<GID>40</GID>
<name>OUT_2</name></connection>
<connection>
<GID>24</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>70</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-3,7.5,-3,12</points>
<connection>
<GID>41</GID>
<name>OUT</name></connection>
<intersection>7.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-27.5,-32,-27.5,7.5</points>
<intersection>-32 3</intersection>
<intersection>7.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-27.5,7.5,-3,7.5</points>
<intersection>-27.5 1</intersection>
<intersection>-3 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-27.5,-32,-26,-32</points>
<connection>
<GID>19</GID>
<name>ENABLE_0</name></connection>
<intersection>-27.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>71</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>20.5,-58.5,20.5,25</points>
<intersection>-58.5 2</intersection>
<intersection>25 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-12.5,25,20.5,25</points>
<connection>
<GID>25</GID>
<name>OUT_0</name></connection>
<intersection>20.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>14,-58.5,20.5,-58.5</points>
<intersection>14 3</intersection>
<intersection>20.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>14,-59.5,14,-58.5</points>
<connection>
<GID>24</GID>
<name>load</name></connection>
<intersection>-58.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>72</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>20,-39.5,20,26</points>
<intersection>-39.5 2</intersection>
<intersection>26 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-12.5,26,20,26</points>
<connection>
<GID>25</GID>
<name>OUT_1</name></connection>
<intersection>20 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>14,-39.5,20,-39.5</points>
<intersection>14 3</intersection>
<intersection>20 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>14,-40.5,14,-39.5</points>
<connection>
<GID>23</GID>
<name>load</name></connection>
<intersection>-39.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>73</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>19.5,-19,19.5,27</points>
<intersection>-19 2</intersection>
<intersection>27 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-12.5,27,19.5,27</points>
<connection>
<GID>25</GID>
<name>OUT_2</name></connection>
<intersection>19.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>14,-19,19.5,-19</points>
<intersection>14 3</intersection>
<intersection>19.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>14,-20,14,-19</points>
<connection>
<GID>22</GID>
<name>load</name></connection>
<intersection>-19 2</intersection></vsegment></shape></wire>
<wire>
<ID>74</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>19,1,19,28</points>
<intersection>1 2</intersection>
<intersection>28 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-12.5,28,19,28</points>
<connection>
<GID>25</GID>
<name>OUT_3</name></connection>
<intersection>19 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>14,1,19,1</points>
<intersection>14 3</intersection>
<intersection>19 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>14,0,14,1</points>
<connection>
<GID>60</GID>
<name>load</name></connection>
<intersection>1 2</intersection></vsegment></shape></wire>
<wire>
<ID>75</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>11.5,-75,11.5,-11</points>
<intersection>-75 19</intersection>
<intersection>-70.5 9</intersection>
<intersection>-51.5 7</intersection>
<intersection>-31 4</intersection>
<intersection>-11 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>11.5,-11,14,-11</points>
<connection>
<GID>60</GID>
<name>clock</name></connection>
<intersection>11.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>11.5,-31,14,-31</points>
<connection>
<GID>22</GID>
<name>clock</name></connection>
<intersection>11.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>11.5,-51.5,14,-51.5</points>
<connection>
<GID>23</GID>
<name>clock</name></connection>
<intersection>11.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>11.5,-70.5,14,-70.5</points>
<connection>
<GID>24</GID>
<name>clock</name></connection>
<intersection>11.5 0</intersection></hsegment>
<hsegment>
<ID>19</ID>
<points>-29,-75,11.5,-75</points>
<intersection>-29 30</intersection>
<intersection>-23.5 28</intersection>
<intersection>11.5 0</intersection></hsegment>
<vsegment>
<ID>28</ID>
<points>-23.5,-78.5,-23.5,-75</points>
<connection>
<GID>61</GID>
<name>CLK</name></connection>
<intersection>-75 19</intersection></vsegment>
<vsegment>
<ID>30</ID>
<points>-29,-75,-29,15.5</points>
<intersection>-75 19</intersection>
<intersection>15.5 32</intersection></vsegment>
<hsegment>
<ID>32</ID>
<points>-30.5,15.5,-29,15.5</points>
<connection>
<GID>31</GID>
<name>write_clock</name></connection>
<intersection>-29 30</intersection></hsegment></shape></wire>
<wire>
<ID>76</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>102,-68.5,102,-51.5</points>
<intersection>-68.5 2</intersection>
<intersection>-51.5 3</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>80.5,-68.5,80.5,-67</points>
<connection>
<GID>42</GID>
<name>carry_out</name></connection>
<intersection>-68.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>80.5,-68.5,102,-68.5</points>
<intersection>80.5 1</intersection>
<intersection>102 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>95.5,-51.5,102,-51.5</points>
<connection>
<GID>43</GID>
<name>carry_in</name></connection>
<intersection>102 0</intersection></hsegment></shape></wire>
<wire>
<ID>77</ID>
<shape>
<vsegment>
<ID>3</ID>
<points>76.5,-78,76.5,-40.5</points>
<intersection>-78 6</intersection>
<intersection>-54 5</intersection>
<intersection>-40.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>76.5,-40.5,80.5,-40.5</points>
<connection>
<GID>51</GID>
<name>IN_0</name></connection>
<intersection>76.5 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>76.5,-54,77.5,-54</points>
<connection>
<GID>42</GID>
<name>IN_B_0</name></connection>
<intersection>76.5 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>41,-78,76.5,-78</points>
<intersection>41 9</intersection>
<intersection>76.5 3</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>41,-78,41,-73.5</points>
<connection>
<GID>7</GID>
<name>OUT</name></connection>
<intersection>-78 6</intersection></vsegment></shape></wire>
<wire>
<ID>78</ID>
<shape>
<vsegment>
<ID>3</ID>
<points>75,-68,75,-36</points>
<intersection>-68 14</intersection>
<intersection>-55 13</intersection>
<intersection>-36 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>75,-36,80.5,-36</points>
<connection>
<GID>50</GID>
<name>IN_0</name></connection>
<intersection>75 3</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>75,-55,77.5,-55</points>
<connection>
<GID>42</GID>
<name>IN_B_1</name></connection>
<intersection>75 3</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>41,-68,75,-68</points>
<intersection>41 17</intersection>
<intersection>75 3</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>41,-68,41,-63.5</points>
<connection>
<GID>6</GID>
<name>OUT</name></connection>
<intersection>-68 14</intersection></vsegment></shape></wire>
<wire>
<ID>79</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>73.5,-56,77.5,-56</points>
<connection>
<GID>42</GID>
<name>IN_B_2</name></connection>
<intersection>73.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>73.5,-58,73.5,-31.5</points>
<intersection>-58 6</intersection>
<intersection>-56 1</intersection>
<intersection>-31.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>73.5,-31.5,80.5,-31.5</points>
<connection>
<GID>49</GID>
<name>IN_0</name></connection>
<intersection>73.5 4</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>41,-58,73.5,-58</points>
<intersection>41 9</intersection>
<intersection>73.5 4</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>41,-58,41,-53.5</points>
<connection>
<GID>5</GID>
<name>OUT</name></connection>
<intersection>-58 6</intersection></vsegment></shape></wire>
<wire>
<ID>80</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>72,-57,72,-27</points>
<intersection>-57 1</intersection>
<intersection>-48 4</intersection>
<intersection>-27 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>72,-57,77.5,-57</points>
<connection>
<GID>42</GID>
<name>IN_B_3</name></connection>
<intersection>72 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>72,-27,80.5,-27</points>
<connection>
<GID>48</GID>
<name>IN_0</name></connection>
<intersection>72 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>41,-48,72,-48</points>
<intersection>41 7</intersection>
<intersection>72 0</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>41,-48,41,-43.5</points>
<connection>
<GID>4</GID>
<name>OUT</name></connection>
<intersection>-48 4</intersection></vsegment></shape></wire>
<wire>
<ID>81</ID>
<shape>
<vsegment>
<ID>3</ID>
<points>77,-73.5,77,-42.5</points>
<intersection>-73.5 8</intersection>
<intersection>-61 9</intersection>
<intersection>-42.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>77,-42.5,80.5,-42.5</points>
<connection>
<GID>51</GID>
<name>IN_1</name></connection>
<intersection>77 3</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>51,-73.5,77,-73.5</points>
<connection>
<GID>14</GID>
<name>OUT</name></connection>
<intersection>59 12</intersection>
<intersection>77 3</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>77,-61,77.5,-61</points>
<connection>
<GID>42</GID>
<name>IN_0</name></connection>
<intersection>77 3</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>59,-73.5,59,1</points>
<intersection>-73.5 8</intersection>
<intersection>1 13</intersection></vsegment>
<hsegment>
<ID>13</ID>
<points>59,1,59.5,1</points>
<connection>
<GID>16</GID>
<name>IN_0</name></connection>
<intersection>59 12</intersection></hsegment></shape></wire>
<wire>
<ID>82</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>75.5,-62,75.5,-38</points>
<intersection>-62 1</intersection>
<intersection>-38 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>58.5,-62,77.5,-62</points>
<connection>
<GID>42</GID>
<name>IN_1</name></connection>
<intersection>58.5 7</intersection>
<intersection>75.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>75.5,-38,80.5,-38</points>
<connection>
<GID>50</GID>
<name>IN_1</name></connection>
<intersection>75.5 0</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>58.5,-63.5,58.5,2</points>
<intersection>-63.5 8</intersection>
<intersection>-62 1</intersection>
<intersection>2 11</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>51,-63.5,58.5,-63.5</points>
<connection>
<GID>13</GID>
<name>OUT</name></connection>
<intersection>58.5 7</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>58.5,2,59.5,2</points>
<connection>
<GID>16</GID>
<name>IN_1</name></connection>
<intersection>58.5 7</intersection></hsegment></shape></wire>
<wire>
<ID>83</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>74,-63,74,-33.5</points>
<intersection>-63 4</intersection>
<intersection>-53.5 6</intersection>
<intersection>-33.5 5</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>74,-63,77.5,-63</points>
<connection>
<GID>42</GID>
<name>IN_2</name></connection>
<intersection>74 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>74,-33.5,80.5,-33.5</points>
<connection>
<GID>49</GID>
<name>IN_1</name></connection>
<intersection>74 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>51,-53.5,74,-53.5</points>
<connection>
<GID>12</GID>
<name>OUT</name></connection>
<intersection>58 8</intersection>
<intersection>74 0</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>58,-53.5,58,3</points>
<intersection>-53.5 6</intersection>
<intersection>3 15</intersection></vsegment>
<hsegment>
<ID>15</ID>
<points>58,3,59.5,3</points>
<connection>
<GID>16</GID>
<name>IN_2</name></connection>
<intersection>58 8</intersection></hsegment></shape></wire>
<wire>
<ID>84</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>72.5,-64,72.5,-29</points>
<intersection>-64 1</intersection>
<intersection>-43 7</intersection>
<intersection>-29 6</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>72.5,-64,77.5,-64</points>
<connection>
<GID>42</GID>
<name>IN_3</name></connection>
<intersection>72.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>72.5,-29,80.5,-29</points>
<connection>
<GID>48</GID>
<name>IN_1</name></connection>
<intersection>72.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>51,-43,72.5,-43</points>
<connection>
<GID>11</GID>
<name>OUT</name></connection>
<intersection>57.5 10</intersection>
<intersection>72.5 0</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>57.5,-43,57.5,4</points>
<intersection>-43 7</intersection>
<intersection>4 12</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>57.5,4,59.5,4</points>
<connection>
<GID>16</GID>
<name>IN_3</name></connection>
<intersection>57.5 10</intersection></hsegment></shape></wire>
<wire>
<ID>85</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>70.5,-47,70.5,-22.5</points>
<intersection>-47 1</intersection>
<intersection>-37.5 7</intersection>
<intersection>-22.5 5</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>70.5,-47,93,-47</points>
<intersection>70.5 0</intersection>
<intersection>93 6</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>70.5,-22.5,80.5,-22.5</points>
<connection>
<GID>47</GID>
<name>IN_0</name></connection>
<intersection>70.5 0</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>93,-54.5,93,-47</points>
<intersection>-54.5 11</intersection>
<intersection>-47 1</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>41,-37.5,70.5,-37.5</points>
<intersection>41 10</intersection>
<intersection>70.5 0</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>41,-37.5,41,-33</points>
<connection>
<GID>3</GID>
<name>OUT</name></connection>
<intersection>-37.5 7</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>92.5,-54.5,93,-54.5</points>
<connection>
<GID>43</GID>
<name>IN_B_0</name></connection>
<intersection>93 6</intersection></hsegment></shape></wire>
<wire>
<ID>86</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>69,-48,69,-18</points>
<intersection>-48 1</intersection>
<intersection>-26.5 10</intersection>
<intersection>-18 7</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>69,-48,92.5,-48</points>
<intersection>69 0</intersection>
<intersection>92.5 8</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>69,-18,80.5,-18</points>
<connection>
<GID>46</GID>
<name>IN_0</name></connection>
<intersection>69 0</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>92.5,-55.5,92.5,-48</points>
<connection>
<GID>43</GID>
<name>IN_B_1</name></connection>
<intersection>-48 1</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>41,-26.5,69,-26.5</points>
<intersection>41 13</intersection>
<intersection>69 0</intersection></hsegment>
<vsegment>
<ID>13</ID>
<points>41,-26.5,41,-22</points>
<connection>
<GID>2</GID>
<name>OUT</name></connection>
<intersection>-26.5 10</intersection></vsegment></shape></wire>
<wire>
<ID>87</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>67.5,-49,67.5,-13.5</points>
<intersection>-49 1</intersection>
<intersection>-16 8</intersection>
<intersection>-13.5 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>67.5,-49,92,-49</points>
<intersection>67.5 0</intersection>
<intersection>92 5</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>67.5,-13.5,80.5,-13.5</points>
<connection>
<GID>45</GID>
<name>IN_0</name></connection>
<intersection>67.5 0</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>92,-56.5,92,-49</points>
<intersection>-56.5 12</intersection>
<intersection>-49 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>41,-16,67.5,-16</points>
<intersection>41 11</intersection>
<intersection>67.5 0</intersection></hsegment>
<vsegment>
<ID>11</ID>
<points>41,-16,41,-11</points>
<connection>
<GID>1</GID>
<name>OUT</name></connection>
<intersection>-16 8</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>92,-56.5,92.5,-56.5</points>
<connection>
<GID>43</GID>
<name>IN_B_2</name></connection>
<intersection>92 5</intersection></hsegment></shape></wire>
<wire>
<ID>88</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>66,-50,66,-5.5</points>
<intersection>-50 1</intersection>
<intersection>-9 3</intersection>
<intersection>-5.5 6</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>66,-50,91.5,-50</points>
<intersection>66 0</intersection>
<intersection>91.5 4</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>66,-9,80.5,-9</points>
<connection>
<GID>44</GID>
<name>IN_0</name></connection>
<intersection>66 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>91.5,-57.5,91.5,-50</points>
<intersection>-57.5 5</intersection>
<intersection>-50 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>91.5,-57.5,92.5,-57.5</points>
<connection>
<GID>43</GID>
<name>IN_B_3</name></connection>
<intersection>91.5 4</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>41,-5.5,66,-5.5</points>
<intersection>41 9</intersection>
<intersection>66 0</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>41,-5.5,41,-1</points>
<connection>
<GID>62</GID>
<name>OUT</name></connection>
<intersection>-5.5 6</intersection></vsegment></shape></wire>
<wire>
<ID>89</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>71,-46.5,71,-24.5</points>
<intersection>-46.5 1</intersection>
<intersection>-33 6</intersection>
<intersection>-24.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>71,-46.5,87.5,-46.5</points>
<intersection>71 0</intersection>
<intersection>87.5 4</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>71,-24.5,80.5,-24.5</points>
<connection>
<GID>47</GID>
<name>IN_1</name></connection>
<intersection>71 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>87.5,-61.5,87.5,-46.5</points>
<intersection>-61.5 5</intersection>
<intersection>-46.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>87.5,-61.5,92.5,-61.5</points>
<connection>
<GID>43</GID>
<name>IN_0</name></connection>
<intersection>87.5 4</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>51,-33,71,-33</points>
<connection>
<GID>10</GID>
<name>OUT</name></connection>
<intersection>57 9</intersection>
<intersection>71 0</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>57,-33,57,5</points>
<intersection>-33 6</intersection>
<intersection>5 22</intersection></vsegment>
<hsegment>
<ID>22</ID>
<points>57,5,59.5,5</points>
<connection>
<GID>16</GID>
<name>IN_4</name></connection>
<intersection>57 9</intersection></hsegment></shape></wire>
<wire>
<ID>90</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>69.5,-47.5,69.5,-20</points>
<intersection>-47.5 1</intersection>
<intersection>-22 6</intersection>
<intersection>-20 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>69.5,-47.5,87,-47.5</points>
<intersection>69.5 0</intersection>
<intersection>87 4</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>69.5,-20,80.5,-20</points>
<connection>
<GID>46</GID>
<name>IN_1</name></connection>
<intersection>69.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>87,-62.5,87,-47.5</points>
<intersection>-62.5 5</intersection>
<intersection>-47.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>87,-62.5,92.5,-62.5</points>
<connection>
<GID>43</GID>
<name>IN_1</name></connection>
<intersection>87 4</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>51,-22,69.5,-22</points>
<connection>
<GID>9</GID>
<name>OUT</name></connection>
<intersection>56.5 9</intersection>
<intersection>69.5 0</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>56.5,-22,56.5,6</points>
<intersection>-22 6</intersection>
<intersection>6 25</intersection></vsegment>
<hsegment>
<ID>25</ID>
<points>56.5,6,59.5,6</points>
<connection>
<GID>16</GID>
<name>IN_5</name></connection>
<intersection>56.5 9</intersection></hsegment></shape></wire>
<wire>
<ID>91</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>68,-48.5,68,-11</points>
<intersection>-48.5 1</intersection>
<intersection>-15.5 4</intersection>
<intersection>-11 7</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>68,-48.5,86.5,-48.5</points>
<intersection>68 0</intersection>
<intersection>86.5 5</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>68,-15.5,80.5,-15.5</points>
<connection>
<GID>45</GID>
<name>IN_1</name></connection>
<intersection>68 0</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>86.5,-63.5,86.5,-48.5</points>
<intersection>-63.5 6</intersection>
<intersection>-48.5 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>86.5,-63.5,92.5,-63.5</points>
<connection>
<GID>43</GID>
<name>IN_2</name></connection>
<intersection>86.5 5</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>51,-11,68,-11</points>
<connection>
<GID>8</GID>
<name>OUT</name></connection>
<intersection>56 9</intersection>
<intersection>68 0</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>56,-11,56,7</points>
<intersection>-11 7</intersection>
<intersection>7 10</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>56,7,59.5,7</points>
<connection>
<GID>16</GID>
<name>IN_6</name></connection>
<intersection>56 9</intersection></hsegment></shape></wire>
<wire>
<ID>92</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>66.5,-49.5,66.5,-1</points>
<intersection>-49.5 1</intersection>
<intersection>-11 4</intersection>
<intersection>-1 7</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>66.5,-49.5,86,-49.5</points>
<intersection>66.5 0</intersection>
<intersection>86 5</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>66.5,-11,80.5,-11</points>
<connection>
<GID>44</GID>
<name>IN_1</name></connection>
<intersection>66.5 0</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>86,-64.5,86,-49.5</points>
<intersection>-64.5 6</intersection>
<intersection>-49.5 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>86,-64.5,92.5,-64.5</points>
<connection>
<GID>43</GID>
<name>IN_3</name></connection>
<intersection>86 5</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>51,-1,66.5,-1</points>
<connection>
<GID>15</GID>
<name>OUT</name></connection>
<intersection>55.5 9</intersection>
<intersection>66.5 0</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>55.5,-1,55.5,8</points>
<intersection>-1 7</intersection>
<intersection>8 10</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>55.5,8,59.5,8</points>
<connection>
<GID>16</GID>
<name>IN_7</name></connection>
<intersection>55.5 9</intersection></hsegment></shape></wire>
<wire>
<ID>93</ID>
<shape>
<hsegment>
<ID>17</ID>
<points>-48,32,38,32</points>
<intersection>-48 19</intersection>
<intersection>4.5 22</intersection>
<intersection>6.5 18</intersection>
<intersection>38 21</intersection></hsegment>
<vsegment>
<ID>18</ID>
<points>6.5,32,6.5,33</points>
<connection>
<GID>32</GID>
<name>DATA_OUT_1</name></connection>
<intersection>32 17</intersection></vsegment>
<vsegment>
<ID>19</ID>
<points>-48,11.5,-48,32</points>
<intersection>11.5 20</intersection>
<intersection>32 17</intersection></vsegment>
<hsegment>
<ID>20</ID>
<points>-48,11.5,-40.5,11.5</points>
<connection>
<GID>31</GID>
<name>ADDRESS_1</name></connection>
<intersection>-48 19</intersection></hsegment>
<vsegment>
<ID>21</ID>
<points>38,-68.5,38,32</points>
<connection>
<GID>62</GID>
<name>SEL_1</name></connection>
<connection>
<GID>7</GID>
<name>SEL_1</name></connection>
<connection>
<GID>6</GID>
<name>SEL_1</name></connection>
<connection>
<GID>5</GID>
<name>SEL_1</name></connection>
<connection>
<GID>4</GID>
<name>SEL_1</name></connection>
<connection>
<GID>3</GID>
<name>SEL_1</name></connection>
<connection>
<GID>2</GID>
<name>SEL_1</name></connection>
<connection>
<GID>1</GID>
<name>SEL_1</name></connection>
<intersection>32 17</intersection></vsegment>
<vsegment>
<ID>22</ID>
<points>4.5,31,4.5,33</points>
<connection>
<GID>32</GID>
<name>DATA_OUT_3</name></connection>
<intersection>31 25</intersection>
<intersection>32 17</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>48,28.5,48,31</points>
<connection>
<GID>17</GID>
<name>IN_2</name></connection>
<intersection>31 25</intersection></vsegment>
<hsegment>
<ID>25</ID>
<points>-46,31,48,31</points>
<intersection>-46 27</intersection>
<intersection>4.5 22</intersection>
<intersection>48 23</intersection></hsegment>
<vsegment>
<ID>27</ID>
<points>-46,13.5,-46,31</points>
<intersection>13.5 28</intersection>
<intersection>31 25</intersection></vsegment>
<hsegment>
<ID>28</ID>
<points>-46,13.5,-40.5,13.5</points>
<connection>
<GID>31</GID>
<name>ADDRESS_3</name></connection>
<intersection>-46 27</intersection></hsegment></shape></wire>
<wire>
<ID>94</ID>
<shape>
<hsegment>
<ID>17</ID>
<points>-49,32.5,39,32.5</points>
<intersection>-49 19</intersection>
<intersection>7.5 18</intersection>
<intersection>39 22</intersection></hsegment>
<vsegment>
<ID>18</ID>
<points>7.5,32.5,7.5,33</points>
<connection>
<GID>32</GID>
<name>DATA_OUT_0</name></connection>
<intersection>32.5 17</intersection></vsegment>
<vsegment>
<ID>19</ID>
<points>-49,10.5,-49,32.5</points>
<intersection>10.5 20</intersection>
<intersection>32.5 17</intersection></vsegment>
<hsegment>
<ID>20</ID>
<points>-49,10.5,-40.5,10.5</points>
<connection>
<GID>31</GID>
<name>ADDRESS_0</name></connection>
<intersection>-49 19</intersection></hsegment>
<vsegment>
<ID>22</ID>
<points>39,-68.5,39,32.5</points>
<connection>
<GID>62</GID>
<name>SEL_0</name></connection>
<connection>
<GID>7</GID>
<name>SEL_0</name></connection>
<connection>
<GID>6</GID>
<name>SEL_0</name></connection>
<connection>
<GID>5</GID>
<name>SEL_0</name></connection>
<connection>
<GID>4</GID>
<name>SEL_0</name></connection>
<connection>
<GID>3</GID>
<name>SEL_0</name></connection>
<connection>
<GID>2</GID>
<name>SEL_0</name></connection>
<connection>
<GID>1</GID>
<name>SEL_0</name></connection>
<intersection>32.5 17</intersection></vsegment></shape></wire>
<wire>
<ID>95</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>95,-13.5,95,-10</points>
<intersection>-13.5 1</intersection>
<intersection>-10 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>95,-13.5,100,-13.5</points>
<connection>
<GID>52</GID>
<name>IN_1</name></connection>
<intersection>95 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>86.5,-10,95,-10</points>
<connection>
<GID>44</GID>
<name>OUT</name></connection>
<intersection>95 0</intersection></hsegment></shape></wire>
<wire>
<ID>96</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>95,-18,95,-14.5</points>
<intersection>-18 1</intersection>
<intersection>-14.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>95,-18,100,-18</points>
<connection>
<GID>53</GID>
<name>IN_1</name></connection>
<intersection>95 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>86.5,-14.5,95,-14.5</points>
<connection>
<GID>45</GID>
<name>OUT</name></connection>
<intersection>95 0</intersection></hsegment></shape></wire>
<wire>
<ID>97</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>95,-22.5,95,-19</points>
<intersection>-22.5 1</intersection>
<intersection>-19 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>95,-22.5,100,-22.5</points>
<connection>
<GID>57</GID>
<name>IN_1</name></connection>
<intersection>95 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>86.5,-19,95,-19</points>
<connection>
<GID>46</GID>
<name>OUT</name></connection>
<intersection>95 0</intersection></hsegment></shape></wire>
<wire>
<ID>98</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>95,-27,95,-23.5</points>
<intersection>-27 1</intersection>
<intersection>-23.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>95,-27,100,-27</points>
<connection>
<GID>56</GID>
<name>IN_1</name></connection>
<intersection>95 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>86.5,-23.5,95,-23.5</points>
<connection>
<GID>47</GID>
<name>OUT</name></connection>
<intersection>95 0</intersection></hsegment></shape></wire>
<wire>
<ID>99</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>95,-31.5,95,-28</points>
<intersection>-31.5 1</intersection>
<intersection>-28 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>95,-31.5,100,-31.5</points>
<connection>
<GID>54</GID>
<name>IN_1</name></connection>
<intersection>95 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>86.5,-28,95,-28</points>
<connection>
<GID>48</GID>
<name>OUT</name></connection>
<intersection>95 0</intersection></hsegment></shape></wire>
<wire>
<ID>100</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>95,-36,95,-32.5</points>
<intersection>-36 1</intersection>
<intersection>-32.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>95,-36,100,-36</points>
<connection>
<GID>55</GID>
<name>IN_1</name></connection>
<intersection>95 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>86.5,-32.5,95,-32.5</points>
<connection>
<GID>49</GID>
<name>OUT</name></connection>
<intersection>95 0</intersection></hsegment></shape></wire>
<wire>
<ID>101</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>95,-40.5,95,-37</points>
<intersection>-40.5 1</intersection>
<intersection>-37 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>95,-40.5,100,-40.5</points>
<connection>
<GID>59</GID>
<name>IN_1</name></connection>
<intersection>95 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>86.5,-37,95,-37</points>
<connection>
<GID>50</GID>
<name>OUT</name></connection>
<intersection>95 0</intersection></hsegment></shape></wire>
<wire>
<ID>102</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>95,-45,95,-41.5</points>
<intersection>-45 1</intersection>
<intersection>-41.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>95,-45,100,-45</points>
<connection>
<GID>58</GID>
<name>IN_1</name></connection>
<intersection>95 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>86.5,-41.5,95,-41.5</points>
<connection>
<GID>51</GID>
<name>OUT</name></connection>
<intersection>95 0</intersection></hsegment></shape></wire>
<wire>
<ID>103</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>-33,-82,104.5,-82</points>
<intersection>-33 27</intersection>
<intersection>104.5 28</intersection></hsegment>
<vsegment>
<ID>27</ID>
<points>-33,-82,-33,-40.5</points>
<intersection>-82 2</intersection>
<intersection>-40.5 31</intersection></vsegment>
<vsegment>
<ID>28</ID>
<points>104.5,-82,104.5,-46</points>
<intersection>-82 2</intersection>
<intersection>-46 32</intersection></vsegment>
<hsegment>
<ID>31</ID>
<points>-33,-40.5,-28,-40.5</points>
<connection>
<GID>19</GID>
<name>IN_0</name></connection>
<intersection>-33 27</intersection></hsegment>
<hsegment>
<ID>32</ID>
<points>104,-46,104.5,-46</points>
<connection>
<GID>58</GID>
<name>OUT</name></connection>
<intersection>104.5 28</intersection></hsegment></shape></wire>
<wire>
<ID>104</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>88.5,-57.5,88.5,-47</points>
<intersection>-57.5 2</intersection>
<intersection>-47 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>88.5,-47,100,-47</points>
<connection>
<GID>58</GID>
<name>IN_0</name></connection>
<intersection>88.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>85.5,-57.5,88.5,-57.5</points>
<connection>
<GID>42</GID>
<name>OUT_0</name></connection>
<intersection>88.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>105</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>89,-58.5,89,-42.5</points>
<intersection>-58.5 2</intersection>
<intersection>-42.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>89,-42.5,100,-42.5</points>
<connection>
<GID>59</GID>
<name>IN_0</name></connection>
<intersection>89 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>85.5,-58.5,89,-58.5</points>
<connection>
<GID>42</GID>
<name>OUT_1</name></connection>
<intersection>89 0</intersection></hsegment></shape></wire>
<wire>
<ID>106</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>89.5,-59.5,89.5,-38</points>
<intersection>-59.5 2</intersection>
<intersection>-38 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>89.5,-38,100,-38</points>
<connection>
<GID>55</GID>
<name>IN_0</name></connection>
<intersection>89.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>85.5,-59.5,89.5,-59.5</points>
<connection>
<GID>42</GID>
<name>OUT_2</name></connection>
<intersection>89.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>107</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>90,-60.5,90,-33.5</points>
<intersection>-60.5 2</intersection>
<intersection>-33.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>90,-33.5,100,-33.5</points>
<connection>
<GID>54</GID>
<name>IN_0</name></connection>
<intersection>90 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>85.5,-60.5,90,-60.5</points>
<connection>
<GID>42</GID>
<name>OUT_3</name></connection>
<intersection>90 0</intersection></hsegment></shape></wire>
<wire>
<ID>108</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>99,-58,99,-29</points>
<intersection>-58 3</intersection>
<intersection>-29 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>99,-29,100,-29</points>
<connection>
<GID>56</GID>
<name>IN_0</name></connection>
<intersection>99 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>99,-58,100.5,-58</points>
<connection>
<GID>43</GID>
<name>OUT_0</name></connection>
<intersection>99 0</intersection></hsegment></shape></wire>
<wire>
<ID>109</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>98,-59,98,-24.5</points>
<intersection>-59 2</intersection>
<intersection>-24.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>98,-24.5,100,-24.5</points>
<connection>
<GID>57</GID>
<name>IN_0</name></connection>
<intersection>98 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>98,-59,100.5,-59</points>
<connection>
<GID>43</GID>
<name>OUT_1</name></connection>
<intersection>98 0</intersection></hsegment></shape></wire>
<wire>
<ID>110</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>97,-60,97,-20</points>
<intersection>-60 2</intersection>
<intersection>-20 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>97,-20,100,-20</points>
<connection>
<GID>53</GID>
<name>IN_0</name></connection>
<intersection>97 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>97,-60,100.5,-60</points>
<connection>
<GID>43</GID>
<name>OUT_2</name></connection>
<intersection>97 0</intersection></hsegment></shape></wire>
<wire>
<ID>111</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>96,-61,96,-15.5</points>
<intersection>-61 3</intersection>
<intersection>-15.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>96,-15.5,100,-15.5</points>
<connection>
<GID>52</GID>
<name>IN_0</name></connection>
<intersection>96 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>96,-61,100.5,-61</points>
<connection>
<GID>43</GID>
<name>OUT_3</name></connection>
<intersection>96 0</intersection></hsegment></shape></wire>
<wire>
<ID>112</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>102,-43.5,102,-11.5</points>
<connection>
<GID>59</GID>
<name>SEL_0</name></connection>
<connection>
<GID>58</GID>
<name>SEL_0</name></connection>
<connection>
<GID>57</GID>
<name>SEL_0</name></connection>
<connection>
<GID>56</GID>
<name>SEL_0</name></connection>
<connection>
<GID>55</GID>
<name>SEL_0</name></connection>
<connection>
<GID>54</GID>
<name>SEL_0</name></connection>
<connection>
<GID>53</GID>
<name>SEL_0</name></connection>
<connection>
<GID>52</GID>
<name>SEL_0</name></connection>
<connection>
<GID>30</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>113</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>-5,36.5,-1,36.5</points>
<connection>
<GID>32</GID>
<name>ADDRESS_0</name></connection>
<intersection>-5 31</intersection></hsegment>
<vsegment>
<ID>31</ID>
<points>-5,36.5,-5,37</points>
<connection>
<GID>33</GID>
<name>OUT_0</name></connection>
<intersection>36.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>114</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-4.5,37.5,-1,37.5</points>
<connection>
<GID>32</GID>
<name>ADDRESS_1</name></connection>
<intersection>-4.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-4.5,37.5,-4.5,39</points>
<intersection>37.5 1</intersection>
<intersection>39 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-5,39,-4.5,39</points>
<connection>
<GID>33</GID>
<name>OUT_1</name></connection>
<intersection>-4.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>115</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-4,38.5,-1,38.5</points>
<connection>
<GID>32</GID>
<name>ADDRESS_2</name></connection>
<intersection>-4 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-4,38.5,-4,41</points>
<intersection>38.5 1</intersection>
<intersection>41 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-5,41,-4,41</points>
<connection>
<GID>33</GID>
<name>OUT_2</name></connection>
<intersection>-4 3</intersection></hsegment></shape></wire>
<wire>
<ID>116</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-3.5,39.5,-3.5,43</points>
<intersection>39.5 1</intersection>
<intersection>43 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-3.5,39.5,-1,39.5</points>
<connection>
<GID>32</GID>
<name>ADDRESS_3</name></connection>
<intersection>-3.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-5,43,-3.5,43</points>
<connection>
<GID>33</GID>
<name>OUT_3</name></connection>
<intersection>-3.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>117</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-14.5,46.5,-3,46.5</points>
<intersection>-14.5 3</intersection>
<intersection>-3 4</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-14.5,37,-14.5,46.5</points>
<intersection>37 6</intersection>
<intersection>46.5 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>-3,40.5,-3,46.5</points>
<intersection>40.5 5</intersection>
<intersection>46.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-3,40.5,-1,40.5</points>
<connection>
<GID>32</GID>
<name>ADDRESS_4</name></connection>
<intersection>-3 4</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-17,37,-14.5,37</points>
<connection>
<GID>34</GID>
<name>OUT_0</name></connection>
<intersection>-14.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>118</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-15,47,-2.5,47</points>
<intersection>-15 3</intersection>
<intersection>-2.5 4</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-15,39,-15,47</points>
<intersection>39 6</intersection>
<intersection>47 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>-2.5,41.5,-2.5,47</points>
<intersection>41.5 5</intersection>
<intersection>47 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-2.5,41.5,-1,41.5</points>
<connection>
<GID>32</GID>
<name>ADDRESS_5</name></connection>
<intersection>-2.5 4</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-17,39,-15,39</points>
<connection>
<GID>34</GID>
<name>OUT_1</name></connection>
<intersection>-15 3</intersection></hsegment></shape></wire>
<wire>
<ID>119</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-15.5,47.5,-2,47.5</points>
<intersection>-15.5 3</intersection>
<intersection>-2 4</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-15.5,41,-15.5,47.5</points>
<intersection>41 6</intersection>
<intersection>47.5 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>-2,42.5,-2,47.5</points>
<intersection>42.5 5</intersection>
<intersection>47.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-2,42.5,-1,42.5</points>
<connection>
<GID>32</GID>
<name>ADDRESS_6</name></connection>
<intersection>-2 4</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-17,41,-15.5,41</points>
<connection>
<GID>34</GID>
<name>OUT_2</name></connection>
<intersection>-15.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>120</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-16,48,-1.5,48</points>
<intersection>-16 3</intersection>
<intersection>-1.5 4</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-16,43,-16,48</points>
<intersection>43 11</intersection>
<intersection>48 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>-1.5,43.5,-1.5,48</points>
<intersection>43.5 12</intersection>
<intersection>48 1</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>-17,43,-16,43</points>
<connection>
<GID>34</GID>
<name>OUT_3</name></connection>
<intersection>-16 3</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>-1.5,43.5,-1,43.5</points>
<connection>
<GID>32</GID>
<name>ADDRESS_7</name></connection>
<intersection>-1.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>121</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>9,39.5,12.5,39.5</points>
<connection>
<GID>32</GID>
<name>ENABLE_0</name></connection>
<intersection>9 2</intersection>
<intersection>12.5 13</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>9,-60,9,39.5</points>
<intersection>-60 9</intersection>
<intersection>-41 10</intersection>
<intersection>-20.5 11</intersection>
<intersection>-0.5 12</intersection>
<intersection>8.5 5</intersection>
<intersection>39.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-21,8.5,9,8.5</points>
<intersection>-21 6</intersection>
<intersection>9 2</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>-21,8.5,-21,22.5</points>
<intersection>8.5 5</intersection>
<intersection>22.5 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>-21,22.5,-18.5,22.5</points>
<connection>
<GID>27</GID>
<name>ENABLE</name></connection>
<intersection>-21 6</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>5.5,-60,9,-60</points>
<connection>
<GID>40</GID>
<name>ENABLE_0</name></connection>
<intersection>9 2</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>5,-41,9,-41</points>
<connection>
<GID>39</GID>
<name>ENABLE_0</name></connection>
<intersection>9 2</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>5,-20.5,9,-20.5</points>
<connection>
<GID>38</GID>
<name>ENABLE_0</name></connection>
<intersection>9 2</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>5,-0.5,9,-0.5</points>
<connection>
<GID>37</GID>
<name>ENABLE_0</name></connection>
<intersection>9 2</intersection></hsegment>
<vsegment>
<ID>13</ID>
<points>12.5,39.5,12.5,39.5</points>
<connection>
<GID>35</GID>
<name>OUT_0</name></connection>
<intersection>39.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>122</ID>
<shape>
<vsegment>
<ID>1</ID>
<points>1.5,9.5,1.5,33</points>
<connection>
<GID>32</GID>
<name>DATA_OUT_6</name></connection>
<intersection>9.5 9</intersection>
<intersection>29.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-43,29.5,1.5,29.5</points>
<intersection>-43 6</intersection>
<intersection>1.5 1</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>-43,16.5,-43,29.5</points>
<intersection>16.5 8</intersection>
<intersection>29.5 5</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>-43,16.5,-40.5,16.5</points>
<connection>
<GID>31</GID>
<name>ADDRESS_6</name></connection>
<intersection>-43 6</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>-19,9.5,1.5,9.5</points>
<intersection>-19 10</intersection>
<intersection>1.5 1</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>-19,9.5,-19,19.5</points>
<intersection>9.5 9</intersection>
<intersection>19.5 15</intersection></vsegment>
<hsegment>
<ID>15</ID>
<points>-19,19.5,-18.5,19.5</points>
<connection>
<GID>27</GID>
<name>IN_0</name></connection>
<intersection>-19 10</intersection></hsegment></shape></wire>
<wire>
<ID>123</ID>
<shape>
<vsegment>
<ID>1</ID>
<points>0.5,11,0.5,33</points>
<connection>
<GID>32</GID>
<name>DATA_OUT_7</name></connection>
<intersection>11 3</intersection>
<intersection>29 6</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-20,11,0.5,11</points>
<intersection>-20 13</intersection>
<intersection>0.5 1</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-42,29,0.5,29</points>
<intersection>-42 7</intersection>
<intersection>0.5 1</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>-42,17.5,-42,29</points>
<intersection>17.5 9</intersection>
<intersection>29 6</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>-42,17.5,-40.5,17.5</points>
<connection>
<GID>31</GID>
<name>ADDRESS_7</name></connection>
<intersection>-42 7</intersection></hsegment>
<vsegment>
<ID>13</ID>
<points>-20,11,-20,20.5</points>
<intersection>11 3</intersection>
<intersection>20.5 14</intersection></vsegment>
<hsegment>
<ID>14</ID>
<points>-20,20.5,-18.5,20.5</points>
<connection>
<GID>27</GID>
<name>IN_1</name></connection>
<intersection>-20 13</intersection></hsegment></shape></wire>
<wire>
<ID>124</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>2.5,29,2.5,33</points>
<connection>
<GID>32</GID>
<name>DATA_OUT_5</name></connection>
<intersection>29 8</intersection>
<intersection>30 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-44,30,2.5,30</points>
<intersection>-44 5</intersection>
<intersection>-22 2</intersection>
<intersection>2.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-22,26,-22,30</points>
<intersection>26 3</intersection>
<intersection>30 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-22,26,-18.5,26</points>
<connection>
<GID>25</GID>
<name>IN_1</name></connection>
<intersection>-22 2</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>-44,15.5,-44,30</points>
<intersection>15.5 6</intersection>
<intersection>30 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>-44,15.5,-40.5,15.5</points>
<connection>
<GID>31</GID>
<name>ADDRESS_5</name></connection>
<intersection>-44 5</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>2.5,29,42,29</points>
<intersection>2.5 0</intersection>
<intersection>42 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>42,28.5,42,29</points>
<connection>
<GID>20</GID>
<name>IN_2</name></connection>
<intersection>29 8</intersection></vsegment></shape></wire>
<wire>
<ID>125</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>3.5,30,3.5,33</points>
<connection>
<GID>32</GID>
<name>DATA_OUT_4</name></connection>
<intersection>30 8</intersection>
<intersection>30.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-45,30.5,3.5,30.5</points>
<intersection>-45 5</intersection>
<intersection>-23 2</intersection>
<intersection>3.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-23,25,-23,30.5</points>
<intersection>25 3</intersection>
<intersection>30.5 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-23,25,-18.5,25</points>
<connection>
<GID>25</GID>
<name>IN_0</name></connection>
<intersection>-23 2</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>-45,14.5,-45,30.5</points>
<intersection>14.5 6</intersection>
<intersection>30.5 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>-45,14.5,-40.5,14.5</points>
<connection>
<GID>31</GID>
<name>ADDRESS_4</name></connection>
<intersection>-45 5</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>3.5,30,43,30</points>
<intersection>3.5 0</intersection>
<intersection>43 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>43,28.5,43,30</points>
<connection>
<GID>20</GID>
<name>IN_3</name></connection>
<intersection>30 8</intersection></vsegment></shape></wire>
<wire>
<ID>126</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>21.5,2,45,2</points>
<connection>
<GID>62</GID>
<name>IN_3</name></connection>
<connection>
<GID>15</GID>
<name>IN_3</name></connection>
<intersection>21.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>21.5,-2,21.5,2</points>
<intersection>-2 5</intersection>
<intersection>2 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>19,-2,21.5,-2</points>
<connection>
<GID>60</GID>
<name>OUT_7</name></connection>
<intersection>21.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>127</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>23.5,-8,45,-8</points>
<connection>
<GID>8</GID>
<name>IN_3</name></connection>
<connection>
<GID>1</GID>
<name>IN_3</name></connection>
<intersection>23.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>23.5,-8,23.5,-3</points>
<intersection>-8 1</intersection>
<intersection>-3 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>19,-3,23.5,-3</points>
<connection>
<GID>60</GID>
<name>OUT_6</name></connection>
<intersection>23.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>128</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>25,-19,45,-19</points>
<connection>
<GID>9</GID>
<name>IN_3</name></connection>
<connection>
<GID>2</GID>
<name>IN_3</name></connection>
<intersection>25 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>25,-19,25,-4</points>
<intersection>-19 1</intersection>
<intersection>-4 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>19,-4,25,-4</points>
<connection>
<GID>60</GID>
<name>OUT_5</name></connection>
<intersection>25 5</intersection></hsegment></shape></wire>
<wire>
<ID>129</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>26.5,-30,45,-30</points>
<connection>
<GID>10</GID>
<name>IN_3</name></connection>
<connection>
<GID>3</GID>
<name>IN_3</name></connection>
<intersection>26.5 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>26.5,-30,26.5,-5</points>
<intersection>-30 1</intersection>
<intersection>-5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>19,-5,26.5,-5</points>
<connection>
<GID>60</GID>
<name>OUT_4</name></connection>
<intersection>26.5 5</intersection></hsegment></shape></wire>
<wire>
<ID>130</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>27.5,-40,45,-40</points>
<connection>
<GID>11</GID>
<name>IN_3</name></connection>
<intersection>27.5 5</intersection>
<intersection>35 17</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>27.5,-40,27.5,-6</points>
<intersection>-40 1</intersection>
<intersection>-6 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>19,-6,27.5,-6</points>
<connection>
<GID>60</GID>
<name>OUT_3</name></connection>
<intersection>27.5 5</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>35,-40.5,35,-40</points>
<connection>
<GID>4</GID>
<name>IN_3</name></connection>
<intersection>-40 1</intersection></vsegment></shape></wire>
<wire>
<ID>131</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>28.5,-50.5,45,-50.5</points>
<connection>
<GID>12</GID>
<name>IN_3</name></connection>
<connection>
<GID>5</GID>
<name>IN_3</name></connection>
<intersection>28.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>28.5,-50.5,28.5,-7</points>
<intersection>-50.5 1</intersection>
<intersection>-7 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>19,-7,28.5,-7</points>
<connection>
<GID>60</GID>
<name>OUT_2</name></connection>
<intersection>28.5 6</intersection></hsegment></shape></wire>
<wire>
<ID>133</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>22,-70.5,45,-70.5</points>
<connection>
<GID>14</GID>
<name>IN_3</name></connection>
<connection>
<GID>7</GID>
<name>IN_3</name></connection>
<intersection>22 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>22,-70.5,22,-9</points>
<intersection>-70.5 2</intersection>
<intersection>-9 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>19,-9,22,-9</points>
<connection>
<GID>60</GID>
<name>OUT_0</name></connection>
<intersection>19 7</intersection>
<intersection>22 5</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>19,-9,19,-8</points>
<intersection>-9 6</intersection>
<intersection>-8 14</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>30,-60.5,45,-60.5</points>
<connection>
<GID>13</GID>
<name>IN_3</name></connection>
<connection>
<GID>6</GID>
<name>IN_3</name></connection>
<intersection>30 13</intersection></hsegment>
<vsegment>
<ID>13</ID>
<points>30,-60.5,30,-8</points>
<intersection>-60.5 10</intersection>
<intersection>-8 14</intersection></vsegment>
<hsegment>
<ID>14</ID>
<points>19,-8,30,-8</points>
<connection>
<GID>60</GID>
<name>OUT_1</name></connection>
<intersection>19 7</intersection>
<intersection>30 13</intersection></hsegment></shape></wire>
<wire>
<ID>134</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>22,0,45,0</points>
<connection>
<GID>62</GID>
<name>IN_2</name></connection>
<connection>
<GID>15</GID>
<name>IN_2</name></connection>
<intersection>22 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>22,-22,22,0</points>
<intersection>-22 4</intersection>
<intersection>0 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>19,-22,22,-22</points>
<connection>
<GID>22</GID>
<name>OUT_7</name></connection>
<intersection>22 3</intersection></hsegment></shape></wire>
<wire>
<ID>135</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>23.5,-10,45,-10</points>
<connection>
<GID>8</GID>
<name>IN_2</name></connection>
<connection>
<GID>1</GID>
<name>IN_2</name></connection>
<intersection>23.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>23.5,-23,23.5,-10</points>
<intersection>-23 4</intersection>
<intersection>-10 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>19,-23,23.5,-23</points>
<connection>
<GID>22</GID>
<name>OUT_6</name></connection>
<intersection>23.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>136</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>25,-21,45,-21</points>
<connection>
<GID>9</GID>
<name>IN_2</name></connection>
<connection>
<GID>2</GID>
<name>IN_2</name></connection>
<intersection>25 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>25,-24,25,-21</points>
<intersection>-24 4</intersection>
<intersection>-21 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>19,-24,25,-24</points>
<connection>
<GID>22</GID>
<name>OUT_5</name></connection>
<intersection>25 3</intersection></hsegment></shape></wire>
<wire>
<ID>137</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>27,-32,45,-32</points>
<connection>
<GID>10</GID>
<name>IN_2</name></connection>
<connection>
<GID>3</GID>
<name>IN_2</name></connection>
<intersection>27 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>27,-32,27,-25</points>
<intersection>-32 1</intersection>
<intersection>-25 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>19,-25,27,-25</points>
<connection>
<GID>22</GID>
<name>OUT_4</name></connection>
<intersection>27 4</intersection></hsegment></shape></wire>
<wire>
<ID>138</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>28,-42,45,-42</points>
<connection>
<GID>11</GID>
<name>IN_2</name></connection>
<intersection>28 7</intersection>
<intersection>35 19</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>28,-42,28,-26</points>
<intersection>-42 1</intersection>
<intersection>-26 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>19,-26,28,-26</points>
<connection>
<GID>22</GID>
<name>OUT_3</name></connection>
<intersection>28 7</intersection></hsegment>
<vsegment>
<ID>19</ID>
<points>35,-42.5,35,-42</points>
<connection>
<GID>4</GID>
<name>IN_2</name></connection>
<intersection>-42 1</intersection></vsegment></shape></wire>
<wire>
<ID>139</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>29,-52.5,45,-52.5</points>
<connection>
<GID>12</GID>
<name>IN_2</name></connection>
<connection>
<GID>5</GID>
<name>IN_2</name></connection>
<intersection>29 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>29,-52.5,29,-27</points>
<intersection>-52.5 1</intersection>
<intersection>-27 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>19,-27,29,-27</points>
<connection>
<GID>22</GID>
<name>OUT_2</name></connection>
<intersection>29 4</intersection></hsegment></shape></wire>
<wire>
<ID>140</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>31,-62.5,45,-62.5</points>
<connection>
<GID>13</GID>
<name>IN_2</name></connection>
<connection>
<GID>6</GID>
<name>IN_2</name></connection>
<intersection>31 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>31,-62.5,31,-28</points>
<intersection>-62.5 1</intersection>
<intersection>-28 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>19,-28,31,-28</points>
<connection>
<GID>22</GID>
<name>OUT_1</name></connection>
<intersection>31 3</intersection></hsegment></shape></wire>
<wire>
<ID>141</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>21,-72.5,45,-72.5</points>
<connection>
<GID>14</GID>
<name>IN_2</name></connection>
<connection>
<GID>7</GID>
<name>IN_2</name></connection>
<intersection>21 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>21,-72.5,21,-29</points>
<intersection>-72.5 1</intersection>
<intersection>-29 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>19,-29,21,-29</points>
<connection>
<GID>22</GID>
<name>OUT_0</name></connection>
<intersection>21 3</intersection></hsegment></shape></wire>
<wire>
<ID>142</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>22.5,-2,45,-2</points>
<connection>
<GID>62</GID>
<name>IN_1</name></connection>
<connection>
<GID>15</GID>
<name>IN_1</name></connection>
<intersection>22.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>22.5,-42.5,22.5,-2</points>
<intersection>-42.5 5</intersection>
<intersection>-2 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>19,-42.5,22.5,-42.5</points>
<connection>
<GID>23</GID>
<name>OUT_7</name></connection>
<intersection>22.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>143</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>24,-12,45,-12</points>
<connection>
<GID>8</GID>
<name>IN_1</name></connection>
<connection>
<GID>1</GID>
<name>IN_1</name></connection>
<intersection>24 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>24,-43.5,24,-12</points>
<intersection>-43.5 4</intersection>
<intersection>-12 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>19,-43.5,24,-43.5</points>
<connection>
<GID>23</GID>
<name>OUT_6</name></connection>
<intersection>24 3</intersection></hsegment></shape></wire>
<wire>
<ID>144</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>25.5,-23,45,-23</points>
<connection>
<GID>9</GID>
<name>IN_1</name></connection>
<connection>
<GID>2</GID>
<name>IN_1</name></connection>
<intersection>25.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>25.5,-44.5,25.5,-23</points>
<intersection>-44.5 5</intersection>
<intersection>-23 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>19,-44.5,25.5,-44.5</points>
<connection>
<GID>23</GID>
<name>OUT_5</name></connection>
<intersection>25.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>145</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>26.5,-34,45,-34</points>
<connection>
<GID>10</GID>
<name>IN_1</name></connection>
<connection>
<GID>3</GID>
<name>IN_1</name></connection>
<intersection>26.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>26.5,-45.5,26.5,-34</points>
<intersection>-45.5 5</intersection>
<intersection>-34 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>19,-45.5,26.5,-45.5</points>
<connection>
<GID>23</GID>
<name>OUT_4</name></connection>
<intersection>26.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>146</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>27.5,-44,45,-44</points>
<connection>
<GID>11</GID>
<name>IN_1</name></connection>
<intersection>27.5 7</intersection>
<intersection>35 19</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>27.5,-46.5,27.5,-44</points>
<intersection>-46.5 8</intersection>
<intersection>-44 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>19,-46.5,27.5,-46.5</points>
<connection>
<GID>23</GID>
<name>OUT_3</name></connection>
<intersection>27.5 7</intersection></hsegment>
<vsegment>
<ID>19</ID>
<points>35,-44.5,35,-44</points>
<connection>
<GID>4</GID>
<name>IN_1</name></connection>
<intersection>-44 1</intersection></vsegment></shape></wire>
<wire>
<ID>147</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>29.5,-54.5,45,-54.5</points>
<connection>
<GID>12</GID>
<name>IN_1</name></connection>
<connection>
<GID>5</GID>
<name>IN_1</name></connection>
<intersection>29.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>29.5,-54.5,29.5,-47.5</points>
<intersection>-54.5 1</intersection>
<intersection>-47.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>19,-47.5,29.5,-47.5</points>
<connection>
<GID>23</GID>
<name>OUT_2</name></connection>
<intersection>29.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>148</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>32,-64.5,45,-64.5</points>
<connection>
<GID>13</GID>
<name>IN_1</name></connection>
<connection>
<GID>6</GID>
<name>IN_1</name></connection>
<intersection>32 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>32,-64.5,32,-48.5</points>
<intersection>-64.5 1</intersection>
<intersection>-48.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>19,-48.5,32,-48.5</points>
<connection>
<GID>23</GID>
<name>OUT_1</name></connection>
<intersection>32 3</intersection></hsegment></shape></wire>
<wire>
<ID>149</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>20,-74.5,45,-74.5</points>
<connection>
<GID>14</GID>
<name>IN_1</name></connection>
<connection>
<GID>7</GID>
<name>IN_1</name></connection>
<intersection>20 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>20,-74.5,20,-49.5</points>
<intersection>-74.5 1</intersection>
<intersection>-49.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>19,-49.5,20,-49.5</points>
<connection>
<GID>23</GID>
<name>OUT_0</name></connection>
<intersection>20 3</intersection></hsegment></shape></wire>
<wire>
<ID>151</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>5.5,31.5,5.5,33</points>
<connection>
<GID>32</GID>
<name>DATA_OUT_2</name></connection>
<intersection>31.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>49,28.5,49,31.5</points>
<connection>
<GID>17</GID>
<name>IN_3</name></connection>
<intersection>31.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-47,31.5,49,31.5</points>
<intersection>-47 4</intersection>
<intersection>5.5 0</intersection>
<intersection>49 1</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-47,12.5,-47,31.5</points>
<intersection>12.5 5</intersection>
<intersection>31.5 2</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-47,12.5,-40.5,12.5</points>
<connection>
<GID>31</GID>
<name>ADDRESS_2</name></connection>
<intersection>-47 4</intersection></hsegment></shape></wire>
<wire>
<ID>152</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>50.5,26.5,51,26.5</points>
<connection>
<GID>18</GID>
<name>OUT_0</name></connection>
<connection>
<GID>17</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>153</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>48,-68.5,48,24.5</points>
<connection>
<GID>17</GID>
<name>OUT_2</name></connection>
<connection>
<GID>15</GID>
<name>SEL_1</name></connection>
<connection>
<GID>14</GID>
<name>SEL_1</name></connection>
<connection>
<GID>13</GID>
<name>SEL_1</name></connection>
<connection>
<GID>12</GID>
<name>SEL_1</name></connection>
<connection>
<GID>11</GID>
<name>SEL_1</name></connection>
<connection>
<GID>10</GID>
<name>SEL_1</name></connection>
<connection>
<GID>9</GID>
<name>SEL_1</name></connection>
<connection>
<GID>8</GID>
<name>SEL_1</name></connection>
<intersection>18 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>42,18,48,18</points>
<intersection>42 5</intersection>
<intersection>48 0</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>42,18,42,24.5</points>
<connection>
<GID>20</GID>
<name>OUT_2</name></connection>
<intersection>18 4</intersection></vsegment></shape></wire>
<wire>
<ID>154</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>49,-68.5,49,24.5</points>
<connection>
<GID>17</GID>
<name>OUT_3</name></connection>
<connection>
<GID>15</GID>
<name>SEL_0</name></connection>
<connection>
<GID>14</GID>
<name>SEL_0</name></connection>
<connection>
<GID>13</GID>
<name>SEL_0</name></connection>
<connection>
<GID>12</GID>
<name>SEL_0</name></connection>
<connection>
<GID>11</GID>
<name>SEL_0</name></connection>
<connection>
<GID>10</GID>
<name>SEL_0</name></connection>
<connection>
<GID>9</GID>
<name>SEL_0</name></connection>
<connection>
<GID>8</GID>
<name>SEL_0</name></connection>
<intersection>19 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>43,19,49,19</points>
<intersection>43 5</intersection>
<intersection>49 0</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>43,19,43,24.5</points>
<connection>
<GID>20</GID>
<name>OUT_3</name></connection>
<intersection>19 4</intersection></vsegment></shape></wire></page 0>
<page 1>
<PageViewport>0,33.5808,338.954,-133.958</PageViewport></page 1>
<page 2>
<PageViewport>0,33.5808,338.954,-133.958</PageViewport></page 2>
<page 3>
<PageViewport>0,33.5808,338.954,-133.958</PageViewport></page 3>
<page 4>
<PageViewport>0,33.5808,338.954,-133.958</PageViewport></page 4>
<page 5>
<PageViewport>0,33.5808,338.954,-133.958</PageViewport></page 5>
<page 6>
<PageViewport>0,33.5808,338.954,-133.958</PageViewport></page 6>
<page 7>
<PageViewport>0,33.5808,338.954,-133.958</PageViewport></page 7>
<page 8>
<PageViewport>0,33.5808,338.954,-133.958</PageViewport></page 8>
<page 9>
<PageViewport>0,33.5808,338.954,-133.958</PageViewport></page 9></circuit>